�      ��Y��H�.^g����V}�$���m f	���I�YBHm��;@Kkʵ2�}��̺���V!!"��Ç�����g_�q��kZW�����/��G\�u�V���X&�?�����_?���ƨ�ݳ�q.�k�{�މ�������!�1����D���������qj���������?]��º�.�B��>�M;�@g�4�_Q�0̣�䀳Q��������_�pi��w�q�B�y��4����^���_`��U�U�4����T��o�㱈�z������_�
��`�r�zw�BϞg
6M<��m�:���(���A�'����ot����,�9�}w�������-�����\Z��p�e�cᷟ�3<��:��q�~�PZ�q7���O�����F�uW�y}FQd��N�iP�B����K?�7����B�1���/��E~<.c�6����m1�����t˼��9$�~��u��뿻:_�O�M�z
��LS�x����l26�7��-ke�t	c�V|�qC2�A?M���D
�[<Wy9�S�9q�V��5���A!��M|1�)�J}�{��'S?������y+�!��C�q��@�|jt 2�D�!r�4`�-�P=�n�O)�s�<@�c�3�S�wsPTg�`'V��Nf�NYL6�A�(dgR�4R�̗!Wv�2x�y��|<��u�d��eF��E�����M8��7����%�G�R�)Uk�4_+�X����V�)��D1�N�����9V��ɖ�y"[\�#A:E<9��m�����0���n�4׉����c��m,I�v�@�rf%��$�#�oD���˚ZXd���sE1������"ӭA�R��H�����uP�`��>�!��ڙ	��Ξ���iK9� � f�+��ʌ��LR�V`�w� ���E�
h�]�vʨ>��.�Ip��	9�qy�Ȃbj�y����+8��t"�a"C%V:���;�̏'/�v_���OH��	�J�"ȟ ����xU�#op'~��	��J��x���Y#h7��58g�@�F���i�����Ǽ\����5�=C�R�.�-f�7|��y��g]�o���{���ϼ�зv�$�����&�N'�/r��ށ~�z��d�E>��-'�'Y�e�"6m������'*�Y��J9(�|w?�t���}��Ȓ��@V<�f�v�A9{(~���xd��l��}�]���8�1���ч�]�������z�ޛu"�^��1�T��Yo�*��"����&y4˃��PyC��d�L��3�� �mf� ��=X��L�^�`�n@a՘ڋ7���șv�e;�����v�UK��0��[8։�� }�9�5������{4Л��2���ʑ�~�Ժ@C�w��M���_�ov�{���.*��I
���J	�y�_����4o�'��A��؃ E�P��z��!��{�EL,,r��@��S{+�6fOk־���������l�dXͻ�^���/KL�<�y��2&w��`�����|~��v�ډ`��vX;`7(�^�dk��1�}���)ؼ=���r6�=�	�ݲD�����6#�O4���/�)X�����>�:���xo���2�/����`'��Ļ��F���^�~�݀gs{��T�%թ�n �l�mLka:,M�0r?~�v�����r��;<���rgz����Bm�֬`-')))�z�w��~7�"��e�%��n��+?Y����Lr��'[8቉>�.��a�������-������'�i��>v���<њ|��`����u'߅�צ/�m^���|o��Sm�nC�2l?m�O���:e��2����[���YO;e����!O�i���v❮�u�Q߱15�� %��5�q��Z,g{l�2�@s��߭ʾz���옒�6�8�ض'��n����$V:�@5�y��v|���z��]��&߁�e�.�]����}(��!'�o�M�C��m�tsko�X��^��)t╒�`M����.~��wt�g�7�]E��رg{�t�/���>,��w���zP/��!# ����b�rgN2b�w!��%���oY�x��χet���� �%�6�uӚDG�����/�}�@��&K���)�]�����܌ipLI� ���8�%�KA/���<��'~���8����@�N��.����偽t���8�a^��^�:�g���|��2�(X�N1>�ys�X��L>��LtM��.�Y>C�����Lr|��ńo^�M�N����b �~%��~:1�MRD<7�.�Iv��
�Pg=���ǜ'���|����>^#>�s�_�3+������dg��O��h�3^���#f��@N=L�|*�
�����+>z����㣩��b���h��; z�8J��~�IV�I6���l<�~���c'�~�5� ?r*����B�{@N 6 ��.�8��|d����t~:�ׂ��ׂ�|�(�
�8z<��C�^��Q��
��騚�|���y=w�q_�{�0�ɉG�� m	�T�,m���b���g;�y��X�������6`���ٿ瀮d�~�����<����y�sy��B#�r-���U��f��b>�9�ǩ����A�<>hy�s�>>�̼r=�k>� ^�ハ�qn���|�~�7�k:7�kwn�����H� j�u�x6}��i^�=���q�Uy�l:�/�2��Ǻ��x>μ��|��Zk5��u�i���Aۣ����4���śl=��h3�^LG�a>�s��M���s���s[Ka�G�G?�<������I^���x3��ƛ����y���|���y^��4��\ϟ/��c>3�^d�q����L��χ��|����/떽��c~������8��A��<i}�?r����=����̿w�;��%�x��絓���q�h;���u�1�5���G��63� ��m�C?_l�?�y<�����^�����6���㷙���3���{go�ɧ�>�������m�k�n�&��_�gn7N�+�s��@���2o�������6������lc��8�>�Z���g淚7��Ӧ?x�n��?z����͞=�ͯ��}M�~���qn3�
�b�/{=��f9}��fsf�|���o3���c�u}�9��ś�=������?�=h}�O��ek�s��)�g�݄���y��8|�s��uÔ||��ǟ2�k�
^�}�㾮 Џ)'�r�/�*�t~����2>�	��kF������I���}�%�?���mA��r=�8��O��������荖K�?�Ku�9/�՟�����ٗ-�y�?��ڜn=�^���}`�����>dt�K�LL���[z>��kPX ����f~cq�;��,��:�2��"g�h�3?u��ρ#877��53�|���z9����<��������53�E��kݣ�[�i�?�����߿���>��3?��O41�4~�i��:���<��g�q��~_�6�������������~�ؿ����{���l�߁������__��r�z'h���������r��S�yw����ϩ�j��x�Ń��ο�3������K���oh�2�o�y��������C���{�����=�����o��N?>�}���|���=m��x���~�k����Z����Ͽ?��UG>���hP��~�"������x�����_����O�2~��ֿI.�m�&/�_ٗ7���c_&�x����=��������mſ���d�_��o�����~`�7�o�ߣ�`��mx���˫/���Ą�����y���̼`^�a���7��L�������� �o����g�3c��c��:�)3��;=��~�\�ݿ?���[3�y� ��x���cO<��$���LO���;>�{�>�{~��s������i}G�L�6���O�M'ٗ8�k�g>L�ٞ}����om�[���?b����C��q�x�q��V<������CM�K�Om��<�f�h����~?�O߿�+^������G���B�nͶo����^�����r�������>�������˺�x���}X�m�<��&�e����|�������O��/}��ㅟ3/>���0���^�������/�g�x����G��>i{��lמ��G�7�>��~�?m ��߭7>���,�?��:>��\?�OX`|�N3�����B�/>����~����Yֿ��%{�텟^��k����|�Υгyڊ7�-����>�����0/�9��M��O��_酟�0����
������|�ӏ��s_��|�_�?�������/�٫��u�m/����x�χMP���v��N�y��7�������_����࿱��������&���&��We>���x���?��A&&[�$���{�_%������<����&��׫L[ޓ�/�������3_�2�i<�om���������h�sb����n����'���3{ɗ�������~ч����=a�^f���}�{_a�_���{����ɯ�?�+���om�g<�F�[��{�
���M.}}A�7�ĕO>�#VH��w��7���ft�� ��9�(�>��{�:��n�
���O����y�g�W�����_��C>�����Y.����WdN��?��/��-w��g3�~�+�'�����������9��|�Ƕ��W�����Ϳ�O}x�Ϳ¿c�_�o��]������ݼو��������ް�+?��g}��-_?�	�{���ׯ9�w~������O�
�����؊_��7>��ͱ���|����c�����Ӌ����O��4k�2�G_�ߧ/}�K����7fy���G<O^|�_��I۟l�K<��u/r�g���/<x��g}�|�=n�N>���x�{�O?����O�>��1/��}����o����:_�[�q��X�������=�}�Ǿ�C|��=y���G��~�m~e_دhS>�����ο�!�
�x���ѿ�L����o��ٷ���?x��C|���B�^y����O|���{���x0��M�� }ܷ�7����|�l+��1������;���9�����X�=�������>�������&7����ٞ}m3>����g-����w�w�߷��:���gOھ�u>��^�}س���b�O�����a�G��w��/��;>�޿?��s��c`�/�����/r��|�k}컘�C��|�kN���{���'�a�_}�W�i�oڿ�!��'��9>�����=�������~�O�a��ϧ~Y���g�;��y�����g�O�5����y��^�+����>�y�_��ٌG~~�����������&���}���ox�#ml�+??�����`Ϳ��!?���|͋_��|��}��.�2񕏛t�O�9�.���x❾�7��W�k��o�b^�U�{������u�?��w1�W9������ޏ��\����/��Wu��Vp������ɾ�����:������������|a+>� ~���;��K}�Oy�'�ox�:ܗ5�������}��s��\|�C|��ȿ��o��/9���/�pOY�
��ʋ_s�ٟ�pO����_�!�����7ۊ�s���/�pO_�"�/9�_���o����+�����1��E.~����|�ǵ|��z����C|��}�'>��ķ�����}п/���u�g��������{����x��.���x���M�ɇ�����?�c��-?�����O�u��?^�c��!���?���:\�K��x�Ͽ͛=��k��}�������X����:���}�����~����k�'��|�����~_�{�5���UzW��ʗ}Y?�����U}󅟟����C|���*���������H��|�{����;<�9�wx��}�����!���?���s_�W9����/�p���K���<�W���Ǜ���3y���5���:�g�{b���
�n���^�m�S<��<��:������=!�� ���wu���9��7y���g_،_���;~�e�)o����)�]�+���}�+�T��\�{b��|~�o2Տ�Ӟ��o�p���+>�&�W�����'��U�������=e�]>�o�����_����?��_�O��k�I���?�!�A̿�g��ۯ�}�;>���X�{����_������3Ɵ��W��������e������:�W�=}��<�w9���?������7�����~o�~��=����?��>�o1א��C�5?��ý�~�g]��u?�lǾ�c}��x�����>�W�]◽�������S�ڿ_�{�5y�c��!����7���}���W}�}�c>�{���_�W�{�A^���_�����u�<Ǧ�������7����c��C|��~����:��!��������r?�l+��1���������c�� �����ڽ)����'�c�k|�}�����?��>���������?�ƿ����b�_�=�?��>��N��]��N>�a����6�5�}����W1q�Z���Žt�ڳ�������?������7����?��>ݿ����s�x�/�p��b�����½��~��a����:�s��c<�1�W{�������5�����_�����~fK���C|g3��g�}�����e?��pO�����n_�{��?�]�5�~~��Wy�����G|&�u������F��^�?�����w��3��/�p�����+{�v?������c�ݣ�/�#����?� ��G~S���������O|#϶����}�?���&�&��u��㱿��=e����y��w�.���O|����!OȽ߯��:�7{��⇿��}�s��	��^����}�X{��)w�i�*�-����s����pO����N���}�o?��>�'��ǽ᳿��=}٫|>�+��������p����z���p����r��}?�;��n��=�b/�7x��M��A<��}��}�7���~���N?�������x؊o��w9��|�_��^��_���3c~����~�?ي_����i��w9��Ɀ��_�ç�������5n�c��=��%������Z̓�ܟO2+=���s$�܏�E����v?�_�O�|?��~ŏX�%_��l�7Y�:�u^���������0��)�>����)`�?=����nj����f��0�l�O���~��}Ϙ}}^����~�o��=�������m��Ϗ:��~=��,������w���^�}Ļ=��s����3.���3s_��:� ���-�2��w��a��W|��i�[��z���������?��7t��xc)����@><o|�~~��_�3���1�W0?;�����+|���O>�ӿ��������ϱ���^��Ŀ���g+������ݜ�kֻ�C6��O�w���^��{E��S�ǻ�s �E�ҁ�!�w����.J�AG���9D��;����=�q��"y*5�1n��T�W�y�XJu�m�vjW��<�G�Zj�Fsh��wE�Y	�'͓-����@��}ui���i�|�{<��-FF�0�T�o�J��+z��k|� ǽ9�?.W���ש���:��~S�X�o1~�
e��PC�1P�w�ǩA�-G"�. D�W*Y�<������9P�޹9F�x7��s�V���H�n|�F w��Hq�}����2�E����}�l���������`na��	��ڈȋ�-�
�zC�yc9������wmh�vFP�]��ե:��)A�ݥ���1���^T7̹ Ǻz��;t;P���6�Lf�KE�qڑ��q�$|��ݥ��wj�	f0���4�K�p��\lƁ\q��S����b��^n��3�^��*��% ���V�$��+25�Z�2���d{[�`�7ԁ����BT��j�!�|�Kٸ��x�a���b}8��mc�����V=�t�.Mֈ=������gE̸.K�ԋ,�0cM�N\	�Y�)���';�\����d�̟~�F�6y��-{��b}�d2V%ڡ�~4B/��v���X�n�-��H�\�*��[n�w�]�J�1�{�,
ɖ��-����N�l��\V��ݚ'�%��+-j�A�X8������3�[���4�k����V!6ܻ�"!����P0^�Zz �i�����|�ʏ���ćV�T~\Btqo�{�fɒ<�E��g���B�!�</Vs�E 4�e�Ipo]��
��XȫJ�Q'u���1B��<&J��]wZ-�\�����Y�W��*�1A*lp�`<��3�ǥ�:��K+�Mؔ�E���>*aƗ�!gK����`�C���<�U߶vg�f��ݲA(�*ң�'M/@[�!�D{SC�7	��u�lW������B:��麅���J�*5�=�J{���%�Ү��0r*�h{)�өGi��v�v�r���čd��r�5���z;�X�}I��m҃���������;�J�Q�T�gSݮł��xj�3�셿��$n��w\;��n�x�FlE��q�ۻB�0����+�&]�-������ć�]`��.y�֠L�e�m�x���8�}S\u��;��q�Ć�c6�p���1��^�1��;��%�u�!���*/K�W��+
��D��xo}<)w3�1�v�W{������ʌW����qԢc�D$����ޯ+����ʱ;Qj �IK��im��T�\�Y��E)m�ㇺ��.L�+�����^/�&�]������0��k�)�T���A�Ι�1��A2�L}�%�n����8�Bl�˧]-7�].��UoEr�l���v\PwuCq���,ݵ-:.�m[��%#�)Gc�6⯌q�m.�/EQNQ9H=�Q��Н�؋�sm�cm�۩E�u{�f^f�ō�v��+w�aV�Kmbt���yZ�#�t\�tD�ʞux�[/,��#��NY)@���cy/���5w��sG2O�i�W��!�{�;gH{��gyY�aW	�q!^����{;p��Qq}����/ٶ%���j̦&�>pHp��0�]E��#4�lW7;"ΦF ������=�������x�/F.t\��Ͷ���%�U�\�YL�e�bv۲��(aW�9���>H���yM� 5��(���i��fP����G��!������L�����r��ѐ�qa�p�k$�
��|y%O|�B@��5E�I}��pr+:��jԊ�T�fmݖ���o�6D���V�^��
n�I=�<��6�pw&0� �Qd��Bw��W���h����R��%�š{jw�Ԕ^ �R̶K�ԏ�w҈:qa��a%��En�U�V6�oU���[�=6D�V}8�Kځ�b�-��s�<�hr_I(d}Y��f����z9���\]J�R��rT�����A���ũ�FN0�ܰ�@�M��	땍�V]bRm-���gD�����#}�e���]X�Pf��f<�n/��J�K�C��`P�`%�)[)~,қ�5Mz}q,|�|���F�Dg�ng�����s�ć�)�%��N}=9��R���L�����v�pS��)���2��� _��/��U�_�(�U�v��K���u t�CC��|Vdgͯ��Sdt���=�>�{X	Ν�:v(e~?�ԫ+�F�m{W��.�Mh��E��5K�-�nO$3B*�ꎡ�vS�s�c�B�b����j��
z<�LϘ!����������3~���v�M1�'�,k�*�"��P��R�!̥
]o4�Q��֣N���5wţ��mc.K�⅛�ǎ'�����"[m�S��o3�*��6#�֋@�w^�1Wn��ı��˸�wPA���t�L���T���~�J�-��ڷX����z���
^�B0�VQ�.wt���y~��7���ZD�
����p3�@<=l��uIn�sq��T�}�_hGxh�<�{r�c�Ҵ���1 qr;����6�o���ߺ���#�B�M�:J������p��C(-���:�f-l���f2�ԧ��`y߇+6���`�Fvگ6Yݜ�^%VBhNQT���I7/ƾ����B,����Mw#d���!u \�BJSD�w3���]�s�~��K�H�yׯ������[r��#�8a��y�7��V�ݡ�ʅ�Ś�6�&����>
ܖNc�C�¦����Qo�	�l����!���o��Z�U��·�����d9����Dܝ�}h��}�﫭M�;�J�ƞ涋Q��ő���T"w拒��jEc��Fu��o�z��/IɅt[89)�$��a�����e�8[��V�n�=^2�ÆZ1���uc�u�R��|�#��G>���O��'�o�j�m>h`�9�ab�_�'��Ƥ@����\J�3~!Z̵x�Mi�j<����i����ȍc�S��X �3\�P⣎��O�����QzZ�.����	���RXnţ72U~lS�I����7���=�,/V!EEQ��a�:��t%�[�S��5e� ���AՀ����k�	U\��3 �tD%�B����6�j�)�.��Q�/�,1.��\�x&{ �k��m~�B�J�n�Rו�l��a�/t8,r���=��N�/�fS�9��u�{g~)w�g�k�q��XO�����[�A偱՗�_S,s��n���s�.:�nȟ�Y>ϊ� vEgY;�3+0Aݷ�������ȑ4���=��og�tx�&������"ע�B>���=�5���ASWFqٜ�����7 o�q�d<a�@���+�Ţ����n.��LJ��7���4�k�ib�"E�_�6L���i�nc�]51^�����MVE+a
����c����n^{]Bm�<"}��)��4\���]�R,6d�p���=�;PQ���\T,��c�*�@섗X� ����I�W;��Y��L����w�H���������hJMdC�֥���z�DrW�r�r��P�z�u��b\�.4����`��< ��>�!�nV����qD_.������ޱtC
B&C�\#9찬 X#�=��!H�������cT�4������,sx���9ھ"�{rT��o����2Y���oC9l�r��d�%�/�.�qu��a�w��K��c=n�u�_]��Y	���د���xhZj9h8B�rw�.#�F���x�Vk�8��&U���ۑ[�w�j�֝@C�UZ�D�_�VQ�_����7�9_�H�|��ǛJ� �4r4l�p��ZQ�'N�� Q�.{���K�?�i�"oyث4ᱶs=�hl���41fryl�ˣYa;���e+bC��$D����n��x�e�2������6j봲�����9�.A��m��{��x�S��-e#���\ ���Uj�K�F��o/(G��t7�RD���xq�F����v�O(�e&k�,�{��f�YLq��;_��n4�[�=�
7V)G��̣�ȲW������5]�A���m��1{�/W5���a���6C!����*޴sf�~z��K���l�t�0��^��QZ���Po�x_\�f��[1���6��W��d
D����K��ia�p��5F�MG��؝�=Q�~�/��G�溭�A�[k\k���4\¼	�%��(U�>��!�����uXW&�D'-g)E�8�
���:�):�֡�V/Av!g{��5/�u9aJ�̓+�a��2VZV�Z��2�ێ"�����|H�o��m�\k�|#jq��ĥ�N��.O�J�	LQU���v���;\�����Q��#���?b|�]��y6��m,�e�����y����|��α4�7�QK�s2D��  \��9^��"Ur�t8��W�lqx烎��wg!"Ӏ��CDD��?���k���u�<��2}��F��/F��H�Z5�iX5QDUG��엞5�)��
��;#��*d�hx�o�h�������kwqO.��\f�;˜Tč��v�ྴ�qO瑘6$��J<���-/�
��7lnw��������~ԡ�\�u=��D�DD��|��ػ��;��)ȭCcX����r�qҤ<��?x����u�T�:F{|�;����QB�͙�ESQD���Rhɑ`s͎��g�������Rcu>�x�j�NL0�6t�x��=��\��|,�G-ƤS90Gf���_-���W��"N�X�m���(G7��n�5�y����=޻z��(_.�ILg�j�ݩ��҂�Ҫ!�@_4g��@��s/s|��%�'z�A9�Ǔq��z�u��w��Q�@$�rXK�|���P��R��|=1����^�n��^x��7����me�:.4�G�j��H���n���BO�� 6��%7���rC�0;՗�@cWNS"��&Ȗƚj�4�6�GR��!u�ބ��h������݆��ϛ�Þ�c���cucF�q��Np���sl�-"ߓ��E����m�'s���a�����a�D/�pA����`�l_ǽdFXWVd#��*3.WW���[����|��J"�}c�NIU�t�DV�V:�N�"����Y诼bU������\��q�F�5�`W�B�R�֫�	&��s>r��Ml/��"�1��{��%ȅ,7�<�ʢl�IEYכk�|�m�)JV�SF2�oB �wz۪nq�o��F2�0
9�.�cm�y<�DЃ�AHR"uk4E7K^7��c�؛x�R;���x��0�] "������/�.�	wHV���M�Y갃�p-ҡIZa����s�e4��Z`��fq�[Y��q�i�1��5�3� �I��B��\���r�0d1\�m[�{	�/7���Y�ZYk�]{/V�ج��ճ������h���=�M�Hgo�U�&m.���R"�D��s�'���蕦BZrZ)��Uu.�}v�P禄wx8�&k�C+Da�fy9R	i������;e�ZŷPX�ju9���RKn}�� 1`�h]�y�Mq�B�k�]���g��5/t��b$=��z���Y�ۂN�Ϸ	1�Z9�b�1�+����8j[hp�xA�-��Ɉ~�����;[�*�hl��`"�&]��a$ۍ�C-"��a.�%�_����qH�,UXub$r�`'s� ��S�>_,�GҒt�2>�r�ݜ�:qb���rL�Il�+>w��*ڨ��lv�.�͕���b4����$n��*�.Кȣjq�S����ʙ�h_w9�t���.ǔ@}�[�ƻ�.�dey�Չʢ�����a�l��h�c.]�Hy�F}0�=�.�]�������>Ee_\g�@�ȧR�N�r�%�2Ūz��]rL��n�
�&���`�s�aJ��ph7�FM�I/��`����l�����lg�u	���C����\�ӻm��oZik�i�x�U��P�,��Nm�=��I�ִ�l�wG_�m_� ^?6�y�+?����uˊ���R���(���H'�QS�T�� ���~�݌[���k-��#�n��MG�ع���$]"�&�i�@Bt	S;��&� iq8á�YP8�1]�m�b��8�	�o�Mw�ߵ����Vx�Z�b��`�$�e{���QG7�-�C&+�(�=��N8ׁ`�MS8_���C�_oO	��)�\��sѭ(<��j���2���.��S�JZH��x�9�Q�]T⠏fp��&A�f�o�
ݖ��Y�q�Y�:��Y���JW�u#�xF�<)��=�����|R:�ĥ��#�"�r�|@Ć��aw����a��l�-K�lo��u�3r�y���Vt�W4�	*<��`ke���Ā�ZR�n,���7���\_f\��!�\�Q�&�U�䑪�gb���~��sJz�p5V޶�Yd�|V��Ks��kQ�*z�O9�Q;&�;��x�ř2��gW��p��=�컣|��nS���V��G|Ǉ��KrmF�p`v��
�g��N�����)Ia��-S;膞4�Z��Z�A�V�L'�{�Ƨ�H�L�����|,����%};��e)�le��K�����CqLR�L���u#e�0��?�6���(9"BǅxA� �W��a׎�nQ�\�3q���ySFE��)ǫ��S�3[��]ñ���`e0��}I���n����zjV���䳚6��l��D�Z�>��X�R�p,ք��燝�}�uFr8��!����F�(�#e����ף��E���f�'�U�wH�f����p{	�M��SDء>�.��U7�g�\�G���~�lّ��H�E�,
Y1̄��-x����a5�����H]hg����l�ؾƁ)o17h�����i�����*�B�Aб�zt�k��r!�L��V��� 7�:����Gd����6�	g�TwQ��K�YL��im��\<Y�21�;�M����E��py���Yt�W�E���P���y��1�k�BWA���پ�o_��e�zh�ky�1:$�>_n��=��_g�p�i�끝ׯ<�Tm\�d7$c�XX�U�3 ��U�Y��=�-��8���Ϝ��t��Ue�n�C�އ!�ֹ�K�b�1y>t"r!Ŵ<T^A]s<�\���uǶ�	��z�/ �L�5��U��:�
Ǆ@�1b�14��zmTu�����mq�����![k��m��g�����.z�����T\ɥ���)�c��YnO~�/4hO�w˸�oxfnh��(�Q.���\�����Cy3��R�Rʥ}����.˄��r��Q�t����r?�7�����%<�;[nS�t�-��3�J�O�F�Dhዳ������S7�$_(c����*�c��j��;k���x��=��f��Y�]�S$�+B��cDɱ��<P���7�8�����+C�%|�SeU�k{y�W���J{���b��$�GEzsb��"�����ɶ��?�#��+T��R��#��Խҭb�4v���<���[u\w��H�w[�����&����,N~s�� q�X�
�nc�]-(���7#Τ������|�A�wj��{U��ckf�0��r���Î������F
��Sp���Y�z[a����lj�F�X�'�DF���Xs=����V7�3Y���ʻ/=��l ���(Kǭ�5�;���^��gZ䑕:�19t_���
V��Q�q�(�dǍ����yd���jɄ�ݥ>ߋ�Xnl�L3�\sM�����b�׳�^��\"3�(|P�zC��L�!��zkOC���¥���j܄�M罹�m�s�v�!��*����1QVj����y̕UW�:��.�O�l����v>Lp}�Z�Q}�`^�
�0ٯ|z�l�`�6�c0J|��s�����}�Ѫ�_�ˀ\���bU0"��zz���;��+�2�8��	�Lg��V8�.U��HS�h���<��.�EC��a��B dN7s��kt\K5N�}ɈJ��:;��λ#�Ij8n�a���0ׁ8�m|�wB]%�#s/�#�{6��+�j7��9F��`�u	�:�ױ3����d�G������q�,ݸ6x%1�o���ƪ܊ң^�����v�yP�f޹�bXEVc)�bp�%���NU�s�la=���P���K���M�=4W#��Yܵ��zs��n��T&lɼ��Ŝg�{��/�r-!��Ƹq��9\d1Gg�,�@�U~����13�͕!��u�p=F�}�\�n��q�覍њ�VS(ky}CD3J?ۉ�O2�B��~��Ղ!��u]k�74�&�)���Z��#$��ȼG�1�p���Ts/c{}G/|*i�ct�c)ҦFd��m8ZY��rV]|�:/���*V�Z���˭5r�G�t�ʹ��F�U��EA��v�3+�k��l���im\�E.��*/�P����.���Uo�0�]�|��s�m�}jU���������Q閷8�E��fb�Go��b�gr��hq�0Ŀeq�ė�Z�E+{!ɗ��b�x��g:��F X��!�j�z��+��jE��|����B��(�$�>�\�I�̲�z�Nߣc[h{ooQ�e�r���k7>h.Q@ӗG=���툔T��MsW!c���ݺG��-��qM�;���bɠ�
-#�d��M6n���E�:H�GZۖ���S���~zk]�Q��*��62�:=&lS�z��q<ز'�Mǽ�Y����2o���Q�k����y6�5��)���{��s^'��P_�Y�@������F��Ll��Z�N����	��s5��ײ��A4�Ò4y���"_2H"I<�"k1�f�ӎ�Cr��ch���]a�s�Y�޺�0-�0e�rQo�^�Ӹ<��#�!�-��Ti���<��s]�0zi�1ۄ��>���nӖwdN"���^y� 8u ��V<���}�����"��Չ�ϸ�i�H���n=����w�^ mܔ-��~T�0����̟��޼�Em!,9�c���^�i�<�ފt!nH�=�s=�;H7�����oA�!o%2s�(������I2���v���,p��&��hz��3<y?w�}λ=������G�q��	��J�:�D+���;�9:���<AN��eƺ)����ۤ�]f���<�9��.Kz�IF�a;e�#
���.t�/�C�ae����3r�y;�C�R�}����LL��/�g|1�wmm��<�'��<ٺNq�y����ؓp���W&~��[�웋>����?i��#X�G@6���u"�c��5���K_�g�/�!g臝�W��k��*�����fyy�������xƏ���q]���*���gxϟ_<z�
h������� � ��s�4���c���q��T3|YK��#���>YdӚt��|�$G_�0�N?�?��9|G��<��7����X����;����sx���E{�/�u��|�}��Rp1�3����<Ȝ�����q��~�z�f�&����W����;�̇�����CT��8��/�+??��3��g��ί��n��5�^��d7�`w?�I`SI$�m���} �!��N����y�<�J����v'��)��r0=A��-����F�([w���z������F�ٯL�0[��Α�h�~�5@:��"��d�VC�k�I&�3�8�k��Q�S+�6�|��uZ�_���]�^?�]{ڼ����״��ƣ�ءo蚰�,���������uIO7j#@���KV��j
���b�ܶ��B�
����̮�o���38,n�K�A D�mԒht�m?�a��-��kx{��t��l@��T$F�R�LwK<葽2��o�:��"�ܑ�W��Ȟ�S�����꾇��R�'���%�Kb��hk�p�H��V�S���tέ��y�T3��%���1S���F���	w�rY���3|�����uiX8��a�6M��i{+H
ϑ���Kޕ�na�˻m�E�����Q^/0�)�Bjw�Zb���m4�wm�^}FV�w����r��y�ˁ��Q�`�R�f¤�˕��,��궺���`yqV���.+�Kf?ƺy���&�D�9��U��ٟ���FV�Q�|.�s�a-~ܧx�ոZ��c����.��Zߪ����2�t^I'�[��T����߃��Uׇ���{��uk���[�
��5��u��c�`s4��s|�z`�Ug"�-�D���^���I����x���|8��cB���w�d�n�(=-�Z��U�z��3B]Q�y�����\kӌ.�;���슏�6Z��0�ԨՑ8h)!�by>�~?l��`	�^^���\gf�,��dL-���ʦǋp��w�O�l
������F(.��R�Y�\^��%��!i�}��z0>8�>�P���._�7����T�-BL,��}������(���m�'u ����nu<𹷞�#�,I[�2��-�����t��p��w�O�9]l
��Hg[9�u��M{ܪ[m\���Hhw��+�V���p��M�y�]6���W���^�QX$Np�wH�ޟ;gV��1���U�3^R�8�w�®T�G$�-41���c��>��D���d�܄�q�J���q9BւƏ�s�YIU���u��K���t�K>6�9S����w��!��X.����W��.�r�o�
�`t�wv+���2������¥~�F�Q�<� K��cb��kz�,Q%X��߼�ӹ�����v�M�B4���QZ$�nXή��f���ܸ{��L��W*q��kN�p~�:wy4P��2r���A�D�sW�՞�L���f�B��J2�d���FA_�VEOӨ�6-f7���Μt�~��K'Ǜ|��<�D��E���ϛ�fs�au��c*ݧ}W�ޑ�������7`pO�H��8\����UV#�vRC'���c:����>���i��^�s^�]����8�%�,tx��*��Shm'N���	��2�ߏ+F�N�)�+k�Z�j���!q�N��V�#��G��Ea�R�p�Es�wȸ*R�l����v�gLr�j��1�%�Y���,��Fɶ�}���f{-��}�]t�izP�A�����z�������b��2[I�n�֗6゜��|T�V�V�&�V�1ǻn�o�+�`�p�,^]����J�j�j�/RB\o�b��Ͽ�W��|��56y�?`]�{źf������/q�K�+���NY�������M>�C>�����{IW|��Xу��RP_h��n1W�hU^U5#,6�:����k�*-�c��|�Y�"hI/�b�]`UY�w�]�~����9��t��2W�
E���[~�,���Jm\��i����Ez�Y���/�¶���(�q8���h�+�T���-���y�I^;s}s�۲��յ]�c�B��%�V��mu�����Es�(^+kH�3>�6�w�^��1��W�����"�&���&�q��{;b���w�"Kw�^uK�.ar�A�u�ojk�q4���Ʒ����̦�y�(T�a���ίJTSk���&	�#;� W��{��t�Rup���r�&�^+c!��"/��z��Ǖ���U}k�r����}��ZHg�T�Gd�}���]>'�*Q��^�0:��򦕾���Q�J�'E�f��p]㡛���n���%ҔW0Rr}�(��V��ci5J"�Ǿmq�E���d9�3�v$Xao\�2��S�j!u_T(]"������ �:�]�S ���6�s�zs㢨	΀B�$A�I������B:�mܞi7��a�j/PLI���z'kN��2�u����N��H�� �nG ��n4��5�[�-��T��q�dy}m��ʶic��Sڡ�:0�;�ƀ�и��|�������1S���jRT�!��0���/�����������C>��@�7��v�t��OϤ �oF��Ć�&\Ӄ�"��P�<����4��=C�S,�6,�;��mo����ވ�w�f<�t6������,�,.�Lu4p�D<�?{�q���o7Y?x���r��S�ĨVR�ep�:2��������]6sB5��w`���6Ċ�+�1�8���>��t֑�wj���|s���č-X.�U7y�����z+2ڀ�]L:�����H�蠑C��x���p��vO�w(1�Jn��ŮT�Av���l���C��,/�7R�r$P��@�8M��g�v����˙�a]�@۳�Rä���=R�|Ȍ�ʌ�t���bRK���d�����a4���9�{���h-6)���7���>�^�5#Я��3��Xs���|kh}��}���{��c~��=2������e���;�\��u8���tiaI摣�����I���%7���2��of�/-A�{���8�h����z%ˢ{�'�C���z��z����G��� ��I�'zb��@�~�~1�uO���n9��[��N�p���\�Й�� D��=��Y����|����)��+f��L��)��|�����U��X̼~g�*�5|�{��Էk���'^d �?����/�{�v�1��p�k4�n�/`��\���%�'��o���f�y"0 =�ΤƝ�b6âj&�? &�����1���p&p�2~�J���~ʍ�xޓ��d��E�"��S>���پ�X�s-�OFp0��1)����Z�d2�T<����_��Wҗ�6�T�x�.�ė�"�����n�!�ߓ�]�ӟ2�|N����K�NY��~�l�K��k����ߔ�?o���/}�"��}�o���_�#���G}��v̜w���[��>?����Vy���?��~K�+_A���~����������w���U�}>�9�����h�᝼��/�-��C����Wy���Y����_qPF��z�'#��N^��z w��:>���o�: |��ԏ~Ճ�����5�L���l��Ys����<9%��_�U�>����9�u�y���놪ɢ�״@&�o����?����Yk_ج�:�~ǯ��y�W�}�Z�7|%���e����̄_�:ʦ�ɟ��&/r�|��Q��W����}�<����/2��s����Ou*�p.ė����RPzw�Y��j�%y��磆���;�+��+�9��e.��������v�L�R�Sr'���^�a���#�`���I���T�G4�9�<�f8��Y4x�O���!N����s�G����{g��<���"������)[��?!�i�a������*���5��?�����6i�����'����j�O���W���qc�b����y|���:J�i�i]1~�K�(� ���'���o����?0
ÿ�5w7�;(na^w��V�6��y�M���__����nb?�~��e�_._Z�:֯׾���]�m]�~Hx^��������cQ����~�����$�9�.>��������싫v^�� ��u���}��c������_t��Z����?���~=MN��2ɬ��Wt���S��-�]]��&��q�&s;!�4��0n����vhΐ����o&`�Hjl�|MT�/Fp.���M)�����ۘZGno�jX�������é$��]DQ?��(jt�qK�"���&�q�V�{l�ٽFj���F���U!*����<��|�)�ȯ��?�����-�� �1R��8+ݸ��G};�����Q��IoD>���m%���������8�F�wK�����X6����ʪ��T}��Ef��(��H�	A�T��~�hhGP�a��ވ�Mg{nC�ׁ���a���ί�[д�kYWIU.���wݙcR��F���(6��l�ԉ��T�b�!_/�2>���
%б��ώt+��@('V�iBʛ���������������fw_�C�8�%��⾲I�c��
�P�8DѶ����R,1dF�K?��HTV��~;����h�#�4����Y�E|7��.����۪9�Bu4�g����ߗ�i��!��x��q(3�$�ТO��ܶ���a]�~�����/�{�n��&_��?D�?s#��s�0��/��p+�)�8��P�0,�b<V�{�M�û�G痥c�[�bư۶�\�[�Z��PB�)%��z�+'6	wiD�������iyT��~��n��X���\2��C����� � P��Cg���I?]�o�]��8w���10/��^�1`�D���Kf��Ǔ&�j�'Jl����`���;��yk�%���;��2Cg;`�7���EXj��9$�/݌�ѡ}����l�tQ:�ʕ�}����N���"�:>���l���
�wA�VN��u�+ιj�"������<�=�c�qGۭ��vuʥ��7;���af��׵Y��q�"����ec�����%VZf*Rj��)���"���+`�N%�2uDa����B1/������d�+�t��S5�7�KF��ȕ���E��ve��Pm�4�� uӄ	�"�`�R��v�1ntZ�T��1-�a�HO0�MH� ����Py�q�����?0%�{�iW��}UF��؅���u7K9���x3���J�ro� ��p��5(����;�����wѤl~\1��}L���j�mxC��JS�����>b��E.�eu����^I(�3ّ�*Y�h-��f����8���t��G�$�W��1����.{i}��-�Y�;�m�d����X�[��҆�V��u���hZ�r/�M��J��7$K[L��}~��r� G��bĮ�B�H(��BR��w\/%m�ǅx/�d����S��sҎ"
t\ZHܯ͕��,�Gl�BQ�:�n�Z�5N􇵾��q�ĬR5!D��E�>D|:���|�)A������+\NuJKͭ�/q�gBh���D�B6�:u�����1]��(�����TW�P�;�8V����vw+����+�#�JQ�؛ԋ�0�ie0bAB$�ɞN},�]��:b/�F\z��keB�x�'����VI�j}���?(�:,$T�v��!�=�=�u
U} �A���kz�/�ﮣ�\�ӝ��amIm2�K����V�d���t:23��{�Zt��wU�N-"�"�(*�NWEt������[�t�QIb�z����lSA�\u��ӽ�i��w37�{?Y������U��:�V�J�M����5��|X(v���n����M�Y��Σ�rp��2�,�=V �;w�x�RE���f
�_p�lZ����Ś��&�z�(7m���cڶf�\�r����"�=B�ix���;���O�dw�r������珗���Ϯ%��<6&��R�<z�&���q�ƞ�M6�'o_��5�z�k�C&t��m<���9��C��R
@�5m,Z׉
��q�R	zyn�f�~�pd�y� 'n壜R����e&���Ay��	��˙�$�����E���)���V�ސ�	f�9 ��Q7)��'�<�����۸E�����;��W��#��JB���q�%>Ѳ�!SH.ODjMۉ�y�����ü������sC�W���M�-�	1��h�i���-�o��<�pS̩��E���s����H��̛"���;��PD|7�Ϗ���y,�J�Y�|T��M�e+;m�����Lۆ����e�ҕ�����`aS��f|H�e�6���̛o��ϥ&Т@2Gմ ���T�~��,�l�"'����M�r��	�t~�0{�3^6�s0����3{+�~�p�IJR����[���gq�g�����΃��S�a*"��S�;Ӎ{�|f�v;�H�!��ykȦ҇�V�_9*�i�lc�������#�3ɇ�����ү�N���}��GT��mN�rkʤ#ճ�|Ʃ�d��(���{{h�{�ҧN�h�s�?�:y~�w?���h������f�ό~�_�ԑ�S�}�9\�Γ��
���;4�kc&�����u�L7)M6f��Ql�̷N�{6`�j�[�����h���������G����?3�gF����3�f�ό���?3�gF����3�f�ό���?3�gF�����ތ64����w)J�k��;��³j�vo{�i����;~�7���rS{ۉ�|�[]��-��=���@s�L䑢�������X�Y!+�>���Ώ:�������
o8�T��������;�p�p׉��F�ƷJ���#�N�#��v��KS���� &
~��p8-�?L�w�Ƿ�3���F���?��t�3��g�fiu����.���q?�鋌��� �o�s�_��՗ �չ~�Q������:Gi�Ku.��Z`���ό�����̈�Tsc0	E��^���z&��S-���;"���g�|0�Ȱ���<��9,����i���f���/�=���Ξ0��p��#{u�8��t;=�R�=a�<�p|>���ߦ1-`�]��"�p�#�����H��o��>NW�[`�o��d�.�L���;b��m��Q��lzd��&�M�Ыh3cJV���q*�,^��}86���3�u���|���������.����3��-(���_c�w(}C�!&���`F���}<8�/P�g��;Y���~@���G�Z� ��!��N�~���<���� ��!ҫ�6��<8�r6��mt��m���Ǖ���� ���rq����卵�'Vx�c-͘�AhK/>�D"��CŜ[��E1��C���������l��k�]��S��bCJēx�S��\��k���+�1�9��x�f�AM������Hd9K�-M����jm�cd-�}���j&���V�W���aҽ0.?�rz�%�j�?�J����G�F[n�:��3u+�N��<H�,�A#�k�SN��"�#�'rN���+M�q�F}wOic#�j>�"9��559�:��a���jA+7$u����w~_3����lnY���Ɨ�T��<�85V^X�l���T���DgH�B��%�{~�X�֢7?�&�u4�:���6��j��"�	��\�dJ�]��*��ّ2j�E���� o�԰�\8D�*�QC!a���_^��z��vgJ��I�a��*���*�:�f�������2\MENW��`8r�	;[I���!��a>��iMX��;��"M֘W�tڦD���&C5�ޗj�B�u���:�M˧���Ke�����[���F�Ŕc�>Җ5�0#eQ�����l	Re�4*f���F�8|%yن��5:ꔞ*O�S܊�U������.��Y�(��oHtp��ϒő�a�,��={��F��S�oT	��w:�K�$��h�������l�@lLmdF��`BaDb6֪����[�vy=�g?R���BX�H�������`����iS�;���Î�
!;��[qm�źq��\ݗ:��I���%�i�����2�#��&q�W���+h�]�Ѵ�j<:7lѮ�{ビ�u7h(e���a��Gk�������<�ٞb�nP6gxľs���uۅ�~�.���u6�4�Īé��}�^~�����xI���"_2Gl��}vΫ]&c7�X���D�f�9ڒ>����$����`�1���-X.W柸v�X���p��f�H�_n�p��'6��tj��n��as���m�> �K㰸�Ay]b�ý!Q���#k�ͦ6��"ZP�ۭ����i8��츐)���Ⱦ�	,޾Q0�q6�g*?&�d��
��%\�X��$��QV���N�* �엧�#���5��������v���(�<�7�����%9p�M��O畷XbWA��c�ú[ap�s��e��
�0Z^xQ�b*�%nD�1^@�B�jӀ�����w�h@�/�����*�R�����3K��-N�c�ǖ�-ϭ<E�����w��Q�T=�Nt:�N�i� IJ,��;����c�ĝ�{T��E�/���-�8)>9F��^+˺����'�S\���%��̹�Hd:V�P������Vg4�+����|WT���:X��D��їC9rъ�B�(ϿdbJe�R�vv݂f�Z�sŭ�E|��j�-�0#!�a]�i��~����~�vĘ;�QE�A���Vab�ّ�1i�2������_)g2���"�Z�G:'e�BEGg9��r�H)�-.I���k���)w�jw�mA�y����J6�e�����w��O�$�a�Rx-XQ� �f�R�����Yh��^z�h���F3T�����-��J��<~#{�W阨 k�ߤc�X��&?�w阨 v��I�D�����
���>c݇鸏o`F���X
���qX;���5�8!��`PdV�����2&�+T�ېX�9ŵ���`Fl�sr��`k��o�h��<�{�ci���ayZ@�;.�NP{>iv�w��C̵�^lv�����������k>q�p�I9����k�㾶��*3�4/fq����,=D�vdn���)�)�P���"��:;�Q9��d[,<G��~�@R�I�k{;V��&�n��D��,v��-��5����	ʪ�_6Y!.ɴ�ܕc%=�$k�����M/����p]5m����)���J�h�\��p���C{9[#��~�ZҺ"9]㜐�$�t�/;cq��M.��»�2,j��U^��J���ݾx;���,���v�tF��n$���{a3R`:�`��tp�\w����|�����D+�$@fp�1Ëh:�m��WǖL� DY�3춲 ���O�:�+}uau���M`�@R,�ts��6K~���9{q��h��xN�j94�$���(��B�)N���.wt4�a���(�N1q�x�>A���r�๚�B�ԭ*/��#L�VV���(�p=��uu:��f��4>���t��޹��C�	l�4��dW�fg��-M���
F-n."�����Kg�)���/ێd��ׯp&ː�ݍ$$�v�5�TNnwq�]4��������֯w -qgL.��AQ�P\� �c���{�)�)�/5&���lm���l�u��z��̾����_{>�[yX�w��������I�������,&�v��k�Ȭ�dBl�d�^��w�lo~`/�����+2U~�V�C����;-�L���Z�c)f��^IC�:��V7��N�Vx,Pk��k��; U a ��������Df�Cܭ�NI�$𷘳Y�E��6+y\��h�H�%b��?�?��ʹ�mI�@�ɠ�k�X��tI\��6"wa�0[$A�68]�#��������b�F�ꎩ=�O�+�S@ᨙ��纐�d�^�K�^ْ�<�L�?�C9���O/I\�B���	�E�^6�O,�<x�e ����J�D{�x�ejE}�} ���J�+,m�aˊ�n�V]֊�����kQ�$��he��+��ͮ���#��c�V�U�x��K�uo'�&=8Z�``E���.�'	��-q�]���)|�֮`��3^є�wO<�̫�!�rA�0��Q3ݸFZr��0�Y5��Ym���\�)�t"���u� j���z�4���B�Ks�qkW���mGrh���jX��p��V��,�?T\b�f�V�R�V)�F,���<��yJ�>�qi�v:������/�����u��NMi�͂��� S��z�F~���E;s�{O�i�ok����օ|�$���)�
��v�P'X̣��ЊLs޸�v��m�k4ܸ�P|O/�#��[,�n�,�A��k�']��s��+Q������ m�G�4w����ٵ�A4;Β���v��|L�ˑ?��o�$�5��=�Rȷ�,�}M�����Kʞ��=o��g^+������?�����e�y�&}����x��?�䥞w�S���~N/p�~�	xX��w�9z/My�P��{�D��X��--���gD*�6'C��#�9�b$�K��g[�
�Rԅ��E>�4���%���i0P�8h��=���pQ��h��#��怩^�w�p̅��[R�2��[$�ZS*�_�����NZ_$������F4A/C&U��0�� �H}ǟ��E��L���mH��Mޕ&|��6�m�ϯm.��P��C�+�B��)��\l�l�ĩ��؄�z˨����޲Ԉ>o𤀷,-����'�B��F���?`�D��L#bm�5���+���d�_�V��D�H���H�JY�C���i��E{���JĚ�
,U�њq�5$� �(^~ԗ8�x����Ey%ؑ�]��l�T����\�R -����a��
ߜa5i�ʍ�\��u6�y��w/-5i3�g9փd���x��3t<��)�����cqHH�Y�k���;�����*v:%���8X�u}�E�M�嘌��:.-j���\�N[K6`��VR�H)��u#��~@�M#ظQ߶�[���*"�M�i�^hFC���X�ud��Zwm4%��*���)`�-a��p�0����9��{gb�-SG����ع\�V��uS����҅��ȶ�xAe99#��}?�J
�+��1��C���έر�Fu��C7����"R�8���87Z>���Qn_n����F(+mW:
���:>!x���.L6b�[���<.�}�i�U��F�b�|s��v���j׮�jFW(�.IH��u�ݙ�����4:�p��Y����w�5և�
����]�tKNY��X��z[�88�x��W9���y���nDL=(���L�w2���3ޯ�μܽn�
;����N�S�N�b��"֛�	}kKʵB�2��h?��,, i�v�f�P,&}��+~{U��mλ�nJ�K��/#�ʔ�HG���K�,c5s����T�� fĊ�m�ú��FX���v���2�|ţ�fŜ�"��rx�W��j�,��
p����f�ʌ���Jܒts��}� ��+~�ꁺ(�@	_���Lh�фPQP�čG�&�)��v0O��7�?�c���ڹ�WiwI?T�����BN�L�]
���� �-: խE����]D��̖���q��g�K	H���?
F�,o��d���һ*r��?\���Zdq@� W�6�T��6�"$��6l&-YgbHo�Dyܛ�:�������.:�����-�z]����"�\n�M���Q=O��q���QV�;�E��b���?DvݭW��:��F�����c�ܝq���&�Fx�P�Go��!	1�{�����X�bG�]��:�}w���V�Jj���˸���
n j�<}u=+�Ւ�2n� ��15��=�������m�gMNA�~u�CeuYŐӜ�X�1e��$���e��#�`6�ʍ�o��Ϛ�)����-Qr��X3�t���hq���vk�# ��<_Cu�ͥV�bP�Ws�����oX�{'=Bx,���_֨�B!��B�d}�����ex����z8>NϺb��L��sӶ �eH�
/���i}LgI�ni�I� �\ݏ{l��ho�r��}&��z�67*	�hu�l��t�\f��o�*�!*�
y� ���38ه�z�p(8N�:׋��D�q�"��WU��x�XX��`?D�����:�m��2;d�&o�	��P�����񌯏�
���xj`�(��ge���hK�Q�/�ӎ�i�8t��׍߷Xiz�z$�5؈��r<K(f��\�~'�F@�{�1Pt(�$�����GDV���t�F�C����������|�O���m��BI�41��Ka�\j��e���� g��T�j���bH"�O/�����.=�hB\�� � y�;��g7�9ZJ�-�.tyY�M��U�d/�̭����]� ��0fpf+G��UNI��U���֮r%Z��ۈw��q�����َ1���wU�Q����B;�z�bɫ ]v��(�*��c�{%�q*'��bo�w��.�wۧ��=r�;�����$��L��M�P�z+z�Ÿ��z��)�]����$�>��"_/��S����N븫�7��w��4Ҕ}N�]�v���+�^��<�a5]�W��c[~jw_�2���-�R�'���)m��`D�[ݲ�����uJvh�Z�1� {A��D���ʸ���|��Ww����F8X=Ӳ�@�r��Ź6MSX^�:-{�����`��(I: ���:��%9w��	�����>�j=��)aY��<`����)��8����Jl(��M��}��v)UߥZ��?�y�i���9�Zh��z������6��g�+W�,��U(Wbp!w��A��jH�����q�7ݳ�(�J�"����8/���@%b�^-^h��;yS��K�9u�����L����am��x�7���l��:XV\���%�� �q�]�;j�7V-�(��U�|�r@4�o�#Q�6�>�	��3��G��-�����.��܆��]r�F��]�˰s.��]'�f�d[���F�`��M=%xۜJ	�0*f��g���j@Gꢷ�� ��t�/WnAI �k3dӸ)��������M��"�	L�������)J�� �xŲ�Dd;R-�U5:�AL��ϊ6dH\���R�;�?�|m{�I�z�F��Hx�)S܆�n^m#ٴ��n�'��	����d�� Xe%5aB;���Z
���� �lskp6]�od|-Nb���67RK�$�/�Vd�@� ���>�SnMي�Z�jqͬ7�&:S���S�5��P��k�踦��F����]i}�n�仗�o�,��M9��E����.�g/����e�H������]<����������~����_w��3/�n?ںGE�%�	�pf�>L��ۤW�R:<n*qz^�F	9
�wޓ3�:���.k/���egL��}J��!?� �0Wc�����R�q�}��j~�Rc2�o��+\�0��Z]�����.����v+J8�pO&�b�*����'r�2Օ2�P���xp���S�����B{���r����/!�N?��|�nG葘����d�9�b����Nl
�+�?���p�(:�Ig��<)�{�#�fM����ؼP�"+�26�d�����NR6'��d�B[��2z{��.[�gN�z; +����z�٘]=`��&�G���ڈw�l;������L��� ��bK!-5j,�:ϻ	{��X�L1��;Yι ���q���-uJ�R]a;��Vj,�)��̭����s۩
�c9���s��"\�:���4:�v7�mH'gG3}'�ޠm'e8���@��`���5�1֜�-l=�X5\Ʌ�づko'�J�Ѳ5ʽsy}\R�C����|� {��������D���a6������9M���J��g�C�H�ツ�[�*��F�rn��!5T��qa�\9Ϊ��F,e��F�3�#K�2�'m�m�!� �p�ۓN��D`6:2`|�t�f8A�C�5K�bz�<|u6 ����}~=Y|�J�PJ/(
���U��<��i��>�#�X�a���T�іNۖ�،$q��=I�k�jå�e0��ֲ"������V�q����8�cL6���WYyU�t����2�U�v�ь� (��Sը{+��P����R��P����$AԾRϝ��9T�o$]ْ�=3����#� 6{��sZ��:A9�_AJ"�����@+V�8��K�/���he�n�/->�@��e5��N��0�����%����'�M���+
��1B-|Ĺ��u^܇������!����"Y_Jj������x8�V�2��V��辘29'K�'#��S,���J�v�o�k<=���iiu豻^\�V���МĚ��+r�-��Z9������U�u�4�y	�iBh���LQ�$�~�#�B��J��r6,�K��Q�P���<6 ~DHʆ�1@�R�]A�`���&���"H��f���S+��_9��X*�wgf�㊙8�G�h��9w��n��[XA�k�*�Gnc�A�4�'�.�V��*��6�ưrw�Y`�~q�g�W-��!+���~/H@���ݰ8.�vC�-��Ԯx9�GO�՜�ӛ}��f�C�T���:68?(���ʡ��?�v!)�ݖκ6(�]q��t�p�_�y����+34�c� b�:�S���-�DB���|X����ј8��8-�k1�`+*�S�&^��[���vE<S��Vz}kx�2Wp�\.-¢�{��nl�0p�v��� P�p�U_bZ�j�j����?��
������ 7�W��v{�b�&�#��kh���b�F8�p,��Ш<��LU�	��z`1��7��H��M�h�r��n�|����x�,�F�=C1ﱩq$��E���"���e�n��$�����u��F�W�q��� \4�z�dʱK�@r�`P�H�uܡ�G��E�^�i�\q4n�+��Pg ��,�n���f)���[��pv�\�� 谤�Uj7=^7�-ԛ9��U�R�G���U)ċ1=��І2�����`�ܟ�_-����M��G&أIl���a�� =*�A���|��m�~��(�[��ľU/S��%5鎴�؄������Դ��Zm�U���p�k���f�
��h�����\�.�``�e�;������)�*�>��-9��A��y��������3^�:vD�j}&�,�ō�R`�B���_fC�{�ל�j�+�6��v��}�gU�7��	,�Y�<V�)9���O8L����q��d�Q9u��v���x��o�?W2�}Ő��g�y������5�����R��&�˿X��&z������ ��>�Ev�ۃ��eB��y�Fg��- '?U��	���KUP�Uo+��xL�/���/T-�}���rљw��&.��4�[@����,8U�1{���Ҧ����a�?�W�mQ���+h@�&@HA�Bk��יkU�U{�:����o��� ���lN؄�!��y�
���9���n�B�JWmr���jCi��G-f�f�R"r���������?���E��7B�u��}v�
��(��CN��>Z��<[���ȚXyȣ��l	݅9�:[����'t�Y^�H�a�v��>M�vF����K����<��[L-���=
U^�LB�iJ4���R^.��sX2��XdZ��_�˰�Z���4nu3%�o:�[T �4������)�=���UQJ	�r�5����=$������
���,&nV��ΠO���3t�)z��jߢ�2����)2���Y�՘���	J������=�xwTU�ﮬ�5��#9�J������K�(��>�/��,��aSu�b0I��N?w_q��c��]7tA<:q�G1z�ם"�I5��x_��s�e��"���r#�5�������Ev��K����2��J�_S�O��s�0�B�џ��ύ����!�؞~N-�l/��X?��p諱v�1S�y9*�0I����՜�g�c����ڝуw8���16�kq�,C^٘����s��X�4R��If��;>��]Ϩv�\}#7�sjlzO�o�1Ξ��U���*x�Ógb٪��_�n?�AG
��?�΁�
�h_c+�F�&G�2�N BF6�@yT�a*�ѫ��E>l���YS� �3�eڱz��-kz={����`W�'��"�����/��� A�a������3ǭ5���!#l���x��fx���!ヤ����39��;���H^�)��;d���[W#tw1g)vc�5c�N�Ȋ�zv	�
y�a}%�^�e>e��wI�{W�/�~�4��Q0�����9ߜ���f�}��a�YXV  S�Pb��l��z��Iz*Ӓ��Ҽ�P�Z[�'2��� ����*ϡ��ͦV*���X�L�#aۋ�	�����?��ɳ�׬P��p_�S���`��[�E�K�V</O(���>���M�"Wgh�>�S�/�NV[�e�A���� ��k�'�n+�q��r�ӗ=�j
�ͅX�C�va���65��: v�g�'�[Ԉ�?�U<�/����:`���H�e��1�u��,�$�I��'1X�W6����~ܢ?������OO�#�`J8����b?��h�ɺ
�ܗX([6�:�,P~�P:��2��K�7�P�1�����R�_��S���g.�D����7$�b��P�������ʅ�PqH���M�c�w���q!�STE�<�yD㣒ZY��[��H�0@�l�J�I�u�
�ࢣ�k5i8=̪�3�s)�4���b�C&檮g� _�� �;�{�-�:@ɪ�4ɦ��T0Mey�I ���rPynҟ+YͱL[[��M���珑�Jдcz^�r; �Wx�1�["0�>;��W>�Z��ܦ����s�Ϯ*p��=)Ŵ!#{z�j�ё'����QG�B����K'����ɜ̿�A�Y���1+��� ��	v$��}�kV�޶X`�Y���	�����.����W�#+�ל �gNX��e��������iV��r��v�ì�����O���l�?�
�]N���4+�w9��?�Ӭ����U�ì���A�������f�.'������� ����� �R�aV��r�`7��Y���	�f�.'������� �R�6+X�mV��r�?��g�����W����9A��8���۬`ř���;�=����-��5���t������~�s������j������l��)�������\ �6f#� �����	$.H�'�� �g!/�n�'�"*�#�˻������c��� U��x$�R�m&1�2��L9��O�,v�-0
~R�cd2k�o1���8|�_Dp�{� ��XR�3Y�'��R�������R(j���|e��uҡF���v���Mܵ�x<�.{?_�~�Z����;d�G�t�v{;�|ҳ��%�>o�Dn+n����:�>޺fٛ�&�WƳ�-�^�JQѹIe�#�0��Uɖ��hb祐��`��d.�����<i������0�I�9Y��cC_��rk�Әѯ�M�X�N�P�[�RH�[ �.�
�L����4.=��C(��_�w�^v�־Ȁ�X:���MI�^�����G]�5�kGͦ5~F
�u���$�o�0��q���M����B�U�ׇk�{�����9�	 �aZ׺|V4t^��� �u�ۏK��m��@~�h����.I/�6?��q��j�Ʃ�����اۆ�:���m�E�Ȍ쨥|`�[�L�9
�7����C��������1v�+u�&�?գe�� �]�^~��x�����e۬���e���C+7�72O<!�c-ר9b�`}�-�O��&j�'���q���\�GQw|Sc���W�Q	�f\�Ql��-M7��U��T�Q��G�K$,�����9<H�s�)�x"�q�Y��>�al<��N�<�Q
3��.]�8���E�oԑjסx篒Q�a�٢x�������ґ���9�ؙ^V��F��t{�Y �����2��l�1�jDR:[|^�u8&%$YF�c�p��n"��_KE��������#�$��u�Y��^��(B	0U�/z�34n� �ljǹ��iZg�Ȥ
��`9�0�#s�>�e���_��	O8\P��2���~��T��FX���&I� ��y��Y��?��Q5�Q*���8��(��J�e�O�U?��>��q�bX�e{`��U��Xl��y��5��R����z��s,�7B�{t�~N�2�s�ϫx����f�0�c	�zqe&_$�\W9�l��J�7��c�7�L~�2%�6�g��v�B؝�#�6$xN��',l�t���fu���GrN.�h�$a�x��^	��%�P�3#Q8zt�t|>mj�Ul��� vi
�d��Ob��:Y+�	W\��͵�Ӕ1ݷ���.�T�$B6��v�>P��PP�o�*F43�����2"4����7eZ��	<����=�p|�&o��4u7�:`7s��k�i�\�g����32N<2G�p+>�UqA�F(�2�p��dI��X�+����0)�y���2����n>��g�`�~o��L�0%mbeK�śZ<��0q��@A��U9B ��+P�f���	~��+01����S��W nGFFӹ��/�:G(Of��O�b�t2�|Sy��%��F]���I0�����a$D_6� 3v����N�,6�7��Yc��@A=%�ղ��JF�1��R
��%��|7ħzv&�Dlt0K�z�;ܦ����A��1K���أ��"R�0�}�a�� 2��ɪ��#7����8Gw*��`O�g�ਿB��aGUZs0*�=�\	v0��$mƬ�3l�O KA��	u݆��I/s�	�i��b��?��In5��i�F�v0�����O0���nT�5�O�Pj�#̋j^�p쐴��
3��B}�T��覊��v�>A��%k{�*�7ib�i�R�ҙ�#�/Z �\�G����׆�v+6>Ǎ2���W���>Oj��UV@��A�+Pt�B{���O_�w�<��3Uݸ��sxSj�ͯ�i|�s<������45�<��9�V��9{3�q�3x�p��$��ܤ��Ͼw�y`��'�>�j�0ǯ���gx��&�%�r�tn�sb���{��:w�s�A����;����i���K;�7������������
�o����WI�{�����o�����Y��ͷp��ͷ�F�9�o+`�~s4�V�5|o4�V o���|[��7G�m0��ͷ��?~w4�V~����|[���wG�m���ͷ��s4�V~����|[��7G�m���ͷ�s4���7��oT�ߨ��Q����F���j���
IW)�O��G�w�)�>��N$�R��	&�c�����&	��%�a��6N����p��U^�^�/C��X4��a��:��~r�(x�����{z���)�ߧR�g�̼K'��̪��@ST4S�������e"�t۾��@��?o��3��	��`S�"R*��:������\?�T�l�ܔ��J8*[a[��ٮ�,�i�a�Qx�W�&�@�O��)���54a��=W�R��f?�#���c4�l���>J�,l���$
N`����ө�{�Tݔ�.a{�-$���1a)��F���;��h�'&#x�Nj�vY	�#a'��ܳ���b�����"S�"y�2�h��n\_��^M��2z��-o;�[`����vc.�Q~��H�!��Kī2����1R�N@B����,t2�aD��Ў��4�{-PtG2 L V��i��%!�/��0��T2�y�8�b��)&?����l����"2rs�ѝ�-�;�w�������_�����?}�����)�
��׺�[�xl��1B��PqZaa� �+�W+����Ѫ&n����<{MP�O�JG��NhbΧoE����Vy���cU��6���KG^����U��S�+�ˬ{=��i#�#G4y�K�S"1�r'����<>���0�����9z�B�][�YV��Y��zy��>�t�J�d��iʷ�����&݌T��E�]9S�L�^K��
7Fo����� cw��k6��F��$��o�~��L�F��׃�TW�Xk�"4@ߦ��+*�6� �1�o�hT�Mb��>&w��@�����q�j[_���"��]s$�j�edI��sD�V�
����	2��ņ���݂���k�7Q��)�;�wa�?>I7��5�	>Sdx׀�y&�͢
�3l�+�pLք��f�`SN�<�K仆붅*�zKR	d��>��vr��c��ڗt�˾W���g���C�Bt�e�n�<��g�7=����b�,�1R�o���ٴ4��9asWX��YLs�ؾ�u�[�S,���p���M���	��W�ҧ��Q#��q� �~M��}l��f:��i���������ܘ<|®���+�e��	,i��1���F4����J�8���hm�T�{�GN
�\��Z��Ѻ�2`F���F����"i����;(��n��$+o�x��p�l�2L�aUt�"�:>$>�Q�!�|7���� U�[Ĉ�l>4v����<�²ۮ�<����!u��>�F�V���zQ��7Y���T�_�2+�u��q�#�k�;�㍻>�x�a����:�����Z��*f���l�ٛ��4�P�"�@�1��It���-��5���L]�%ڈ�.6u���/�j�����$��b4��Y8�]4KN�o�ie~��+�U� ^��F��򌋏�pQ����t���o�\�|�	��ݲ7�m��4����6��)�U�BД�v=F�9W�T��lB/�s�Nx���=g�H����0V+G�ğ�p��Ǩ������Άg�����(hz��A<�3a��OV��	����S�^�\G��3�F�OM��C�53�܃�W��C=�{�=6�CBOm�4x$&���r�<Tɛ�w�c�<��ɍ6*��2�.���:*�^�����,Si�&w�עuCi����[�ē+u�-�3k34���%[�U���cP\�8��8�S��������SCz��o� ]�/����g���(������́��6B���^ށ|��}�����󙣷�����C�3��/���K-�(ک3�s���N��;ƆXA;?�¬��H��U<џ��9��"�x�/�+������{7��U6�姷��I��֣���g���� X�9ǡ'R��ʉ]I��K	��E۩r*��9"rw�����e!��dKJ �؝³3���"�_x�f_O^i�z������P,4�4�RKR�f�f�su5�̯���Lfb�jwp���c:� �Mx����9\���}�q�'cm�̵֮��Vv"�	Í�r�'33g���c/�p�Y ��.ׄ�%��, W(k��'ј�^Z�("]�X�&&����? /��B����%��l���U�.{_{���(e0v����Vhۃ#R��m�~�=�K�,��se�G�}&S�{��|�ok\q�c��]qbƩ5�OZ������E�F�nC.	%K2�ǒ�%G�Y9�ȼp��M%p���E��v�̛�������\��K&٫h�X�l��B�uO���%�/�^E����Xah3S��P�{.�`Ɓ�V?���mn �6�����ݕX�{i�)��Y�P�Ԭ-��'m�`��i1��n �3�ͷ�8�Q9�/�	_�eܝO���g��;F
-LU��|^���ugq��CǮ⼷T�}��0r��'n[y~x��bx�`�#Z���U}�%R���b��j�~��u����N���4m�Gt�����8h�G�g�tt��R-Mj�E�[W۝�#'I��^���6����#��Ti{�k���z޲��?���skUx]Ti�ӿ��GU��?�g]��?��� ދ��Z�[����������?+ݻ��-K1i�(5�#�R����h�L8:����m��]]dT�����~\��F�ټ�}L�1��@h�V�d�ٵCG�۠r��G�U��]��Z[fo9�l���%c�24��N��U��.�I�C<r�qRT$���	ʻ ��ʴ�����z0/�� �V�xn�f��L���VXpy2}ܮ�Ǽ�- �> ��=bn��C�j6��K�m�)�	S�wD�P��[�����|�mўbgh��j��T��ݜj`�(��JZb䡾�~`F����q����7*�mf<*������ 3x6}��}�ڳ�0	�pL��Y49�2�3(��Fk'Mp��$:"��l���ӥ��ăp��?����¿��Q��#Apa2��*})�V�U����f��>2�,���@�]��־�����f�d���Z��?��$��e�L�	$�g�~��TD���;���243�PK�C�xnHUn.�Гd��=���������&3��+�O�3���Z����0���
���m��Yzn9a�@���u�=,��)��M/`�����@��ͣި�j�=���M�>a�%w]ԥ>Y%cZ��H�⓵8i��I1��R;�J�k��E�,9rfw�H%0mkKΟ��4�ys��e�}�S�|�<��{�$�	/���߱�\�N!lMЧc⑊��w��PƝ��A��w�����|��� u`r��XN����{��/�C���V������u$��������7������'��h�r�r��P���{�߁i���ZW/u��2�Z=@`J1		���/����dȷF5@���C(�-�{��'��"�oe���t]~c�d�R������~ԛ��]W�xGt��^Hܭ�_mZ�$�|Y����-"��<Íxނ%�3%�:fɲD���c�e�b�f�n��pHҹ�y����IS�-�
�� y��R�����fr�y���ߟRؗ��j��	�(V�ǫ������rm�ƀ���1�G��f�f*D+Aέ���a�'��{���G��H�����(�V��9㺷��*[ƸS����=���{���z|W�u�aϑy�#�It��;������>J�ǾK߭�\D��B�$�CvӃe �6�?�����VL� ����c���T4��LV3�2Y���*�/4vkj�����z������]���?Hȁ�T&���x����3�Rv��}۬�c?V�ص������BCD�I���T��K��x~�q��N?�9��<:��r�#��9A�3���i�Z[�xf��E�P/����`7�8.�p��p%����|���J��>�-x�#}�LU
�Y�zF3	�������:��朂IO�F�_�_�:�]&ସ�:��Iݦ��ByK��6��JF��a%�0�1[�8�PQ����=��C�������>8u8$)c�X���7��9`������xq��e���#-��7Ƅ�^�H݌��}��w�o��Y����?8%+�Z-6�����q༁����d�W3��,�
��{���#���o�0���8��h-ʴ��o=>��3f9Ű�!�h`�+�v�j1�N�!��"}�jqFB���¨>am;w;��?|F�o� �ִ��PeX_�9�R��R��mt���Z�[�}��{�%%�-_xG�U�7����^���w%����z��*lE��C���wM�M����j	d9���0>���[��0'sr�&�B���q孼��(q��s�Ll��h�Єj�^n� <��0N �?1]�5/�7�=�f�w�������`�q���ק,y򐎏�OL��{[{k������H�Z��sO��no�>�p5�>�)��N>������� ۵�>�=��F[�|)�0��1ʴ�ic�hdӨ�;�#�� ���>��[]�Li��A�oPf��4W}V�����;�r5KQi�2�W������#kQ�7�R�>\���_O�ۦ�����R�u{���[�[LQ����$� �Eu��������{/ȃ����F^��lTy����y��O���2M슶ȥ���L�{X5����^�y�nE׃]��ұ�F������7�Ѷ�����)I��� 0d3%4� �Q�9� &�hf�-}��}(7N�\�lXmӽ]=�[Y�2�ю&4"i7{ܽ��'�x����-��^����N�[�syrV��Q�73���dA�U����O�M��B����-��sf`D�u�[F��`,7L�,��9��fi���&?��%�t��ߧ�\�i�� �ۮ���d.�Aa�ޓoJ?	�綳�D�3y0�rVY���>�����Xq*5�L�[��YA��{�A��lN6��E�<��h5���Z<��)��`�G�յ��VD��f�����B���AJ�4�d�I?�TpW̶���'\���V�w�}.�s������ľY�-�4�(������X"��MW�@�	��>�.c<�i3��՜'�����|w5�D׾d�{����Ot�f1}�V�3��x�0�'�NԔ�a`���~L��3ϜB���B�����/�*,���Q�o�wĝ�=^o�	���JP> ���B�;��v��S�Q�����A��K�]��7�c9�p�Z1��3��B]�R�tr�w��Ulǥ�0��d�R{�b����*�S��tK�GT/!s&���?��ߣ�6�U���NZk	�=_�rΕ�y�Dm�c����t��/ۯ�U�H�;>[W���< �~�}�uMD��H�=@��m�wb����/���3�R����h��Au֘�C���b��'k���� k�7,�cѓ���Z��ː-�V^�ѭJC�����#���8/dg�x6
@b#�}��yN�ܼC8�����^�%����9�75W�:$�'2E�D��߻[X.�ּ���q?e�$N|��s�+����d2�'d,����L�h;S舑��_�o5�y�|ֻyO�7Ųa��$�\X���!�ϋ�(q���u3�ֻ��ҽ��O��0��]#z�i��w9 *�m.����Mؠ�Q>ϑ�{("'|��|��I���1Fv� ��q�$E?��L_��q��S�w��u�6,�}�i�:�UJ'kF3�ԡQ#<` Θ5�����%��uZ����՚��&�L�+o]�3��jy4w��)��뇨O��[l�!C�Z!��*��$787�vh���7YW�%���)N�����;�w�H(A�d�Ȁ��Fg'!�J���Ӱ��#��O��e��� ���+ox��nX2vٲf�a�#(�.K�C
�p�NK4�Y���c��PP�.�C�����+��/�'`�b��O��瘍���O�X4l�=�FZ\�S	H^�o5���[�;���\�E�G�B�����@�9�%�>֬ʘ�)ƛT�:��!킹y�(���P�Vu����=ix�A�@L�H0�+l�/��,*;LH�܎@���y'�-
",��xi������_�#��kn��Kn�ˆߎ!� ��W�'�}��_k39��;i����Q�	x2�ү'|��{ల�E��8uz�>��b��x���߫�s	t��9�K� D_�IGk7W���*�S|<�,�	��O����Q�>}����׋s,������P�ի��z�\�e��e���4��0X։�Gzdo.����ax�p�/���߸�+��Gm�5k�o{@%)�;rZ�5Y�I���:���{����=�� o��j��}c8U^	�}��g�ٗ��>Dq�tG~v�"Sz�Hv�).>�O0aH^��"��`�<���Gmr�4�T�v�[��`�,�����.	�?>���&��|6_݉��2�]	Pń�Ja/fo����vp&b��&枳�˼���O� ߿g���秏q
�C�8����'\�}������N~7��S���cTC�H�����7�O�_�D���!�@�p6�>c6�ͼ�l�>r�!f�_���pKk݊�,�O�Bb"�R\�V�P7�(�;w��.Z�������b���"N�����	n^�� ;gP;���ݘ�ݹ�\a���d:^d�7t�[����̒�pZ]��Ϳ�j\ܦ^�	!�����S���zp�G�w��[S8#>yQ
>��R9JM��x@�w	���)���5�$��(W�������Q<Gn�8�Q�jE@ĥ��Q�j=���7i��(� �S��<�^eu}DF�D�P_�!�.>3��������,�@�_2�r���{ג��QpC^S��p>�x�1)�PhO~i5Z��j��F��5����]yG ZhA�����(N���X�}ZU}��F��n���*�T>(�B����%)��=ළ[}:\��o��AV�ꆶ�x�A6�T�.6�2��6��xl��b���,_����Q�=u�i�[�{��ϨЖrt�Tጧ�eϙ��t?东V)NT����u+�\� N kt�w~+b�7�hC�B�^jT��bʏ�s�|Q�&�	��;^�F�1 X=E��j�D4⭑}J���#�1?2�z�}<ۚz\ö�oJ��v-eʆ_D�J���8Tؔi�`^�Z��W�p����%���<�l�m��<�N@[�J���$�'����?�6�Bۖ���J1j��_�ʟ�����`�7r�G)�"�da�O�/n{ķC�Ub.����^����y�"�(�U�%<���*H���D�@c��Lhi��u'i͟g�hcO����N�D{���3\m'��B���N��� �9R_k=���b9q\̨	W�D�NƼL`����Q��L�d���7�e����b��r�at��3�#Ҽ u#��!q{�w�4�) �U�M-T���۲��ox����jo>q�_yk	P�Q���,]O�	�*�U2>E%}|�Q2��[�!��+�"RwzǵC:�|K�>���Dk~�{9}�������t�{�Km}<K\�w�M�<߆�QN'�%W���z7�zG��ɉZ=�Jr◇�w���v=��w31�����	�?LC�V�n�ZhG1�oD�W#)����SdG��O@�ؽ{N@�=5R�қq���W�F�[a6>ew1�7��'8|�f����SnĨ8j�`���V�/]��-�72JC�Uf}��~,�V��&T2��u�(����s�cmx<�R��|��gX{��wJ��򽏆�0d[�V��1�K��#����zTC���ݸ�o�#{�̥M���[4�ѴHNq�f�Bv�GX�%��K���͇/��vo��}�j4�\� nXJ>�8f|�4�C:*,�b<��xd�a�-���N�Q�! �j�������U��e��ݦp�ƾέՇp�rV��*́���H,�+jO/�e ��Bo�ꚉ,�o���:֓ibڗn	���m�#ƍ�kS2�Q�3�C���U�w�eߠMSy� �တ>�1�� ���r\�$o92��4/1:��P'�r���O�%�=S`�%v�L^o���ԒR������ƻ�#�r1a�?�b�D�a�҇���j���M_X��\TUN�2����=��g�A�ڽ$�N<η=E�|Ά��<��#�y;�����f�д�w�h�8�X�\�N~�i�����Rh�ǎc����-�i�X��T�b�� ��Ks'��]x�ٕ��5���٦O��~	�����<�V��`����V%��M�a�TzO)�}�
/�d&�szْ���d1�M���o�04�{�dh/�ik0^���`M���s����I���uu�TI�R��x��UE���P�����tDc8��G�0�$ǉ�V�\�x\�œ�:.�Um���+��C!x���:��U�f�W�Qˎ5vN[1���dm�/��űҌ�j�=Q�ί�^Y��=�6����㓷v7�}�(�{8�U(�@-�لM���Entc�4�T�GO���
�ry�^� n_ГR�*ǧ١%��$fR��
���Ŷ�;���		~G�Rn��9F>�Te�A �BWy3~��D]g`������
�6 �J��ը�R��z�,.�9��_^D�7`���39�u.U�;�l�S�'<x3��Sp�V���Ĕ�U4W�0�dK��~+:倪�� aM�~r��HcAKN`0�R^��G��o�P>!}^7�-�\�h�������V���RYJ�,���ZvT}m1C�����3G�X���ǐ>c�y�M�?�_Z?��'=���Ut�{�3��(i�xJT�+�BY��"j��JQC�r��݋�r`�v�� �5�Y��Џ�{�G�w�_���w"�vn�CS�kR�B�A�#���`6�x�[�Ř�f+��CpM�q4�1;��Ȣ����{C&��/�:�Ɠk*Ҧ9B>���V��6�yT^�E��O��#={�,�쫟�#�f�_��g:�� 6>c��X���7��k�%��q�o��2�S�趦k�~R,���x5y��3L~�ey�~��^�Ԗ��3":��fS}R��ߍ58M�fi�|Ȣ,����;��:T�d�=w+�����o�s]'��#�ܢ���<��9it,�F;��;��*�j��~����3��y^��<4ax�WqP�Ad��QZ�c٘#�VNq�p��L�
��-[��Z���k����I̯7;�h�7B���]�}�M�\�����I��`(m�ѷ������G
��F����O�m�<�Oa�j}�lZB>T�	 �?�A#�
�ȯ#��3�]�q��f��ܕ{�tM�:|��ɐLg����0������g��=���%��~+:�i@/�| N����0����qy��X4���������[I������I|�,�5@AOrZl���9;vi�=�`v1}R�y�z��`j�:�����xMxF�/(@�o<4Y�S߻����1��� �'R�~�!m/*�I��&�7y�S��Ų�-���V�o�R�A�"�_�H��~�>��a?�F@l�#�<!m&_6C��u�M��[$M;���WGv^	M�wѮ���OVqs�F�Տ�{%sz��My3�&1�1��n�2�o�u���;���:E풻��a��� 1:�x�[����)9�.�	�Q�7��So��u�s�F��ʮ�Wd�G�d�M8��K����Mj?�*���\���ɝEZ�9�m�Le��*�'�znl���y��U����1��̖�מ�>�BIw��`���N�Lk���[��(���oQ �0�_  �`n"�x� �a�LD�=���:-��Ъ����/��I.�h�_�H�)�X�|��'h���K��!^�$Bh�M�Zҟ�u�F�\��� �4�K <`0�&_Y����JIy��u+�N�]��Q#��; Z�c������DG?�U��o�/83���7�A�:�H��%ep�r�k{�1�#[)d� ��۰�I������fS?X7Թ3{���i����)�
f�&>�}{[Md��!ߡ��tY���s�Ҭ{��h�6`YU���k4�ܞ���d%&T.����Q*9��#k����H�6�UG��
2'���(_3�A�[��+�-���Ϛ4��M5���Ѐʬe�Sv<���;^���G�}�d�W�L!�<�t����d�E�j�}�$�,��>>�A�C��&���X������u��������#��d��AF[=�3JĽ�op�M끚��]��������d���(!�%p���>7�o�Q�!�M	3�q��Rװ���Gv<e�x�-'Utr�g�^�$P��r| ����~��#q��h'VsQ�xE�8Z�w���=��S�׭��NWC�����Q�؆�@)_5TZ����^(O��>����*b�����Heu��9�Γ��MX��/K�*��CZ��e��04vN����X5�%�� �"��=�|�kYi2V��~,D����kڴ�gA�t����c���$G�U�+�����ҝ�#i��Y������Ek�.���8b�>Ip^�!ҚAț�o�A�^k]�6��G�݉U�q���s)�%���g���w��4���a ���X�����Jp,@mq� {��~F�d�Z#Ȍf�L?ٖy ��x�\��+�Z��0�ƲC�{7t{��\&D*���~$�x��II2�~�N`�X�j%�^�H� E�u�)g_k��~��}����ۅ��%ݫ�n�Y3öbV���$���l���
%E�������]A�h�ώ�f����ǭb[�࿒�}�R*2, �v0%h�y����K���c���aK�����Y�H�0)�1�G9_-�O���C0�����K,A�2�T�9ƃK��T��8j��i�[oٽ6��u��&�d^VO1BԔ(�NɆ�܍
8rh9ij�X	xcz�(�y
��a��^��J�#{}�tD[��ERr+�6z��b�3�����jd�w��T��"g���ZkÅlD/'��v�	�g�bz	O/_�:Į���@� ;D��E'8�(���(�u8���-i�����F?�t����<5�FƬ7	Xdʻ��Q⤃����5����ek��"�,t�������
.����iw
@�M�(�Cx��b#�LO�M����}��f򣓌�AQ��5����L[��IC�0�)��W��߼��ݞ��G�d�{�G�(
��ݢbA��cc���M�]��5�8�i���z>�9�EQ�<|�Χ�N�qǎ�CR�C�8і��ݸs�)�т��`�,Ida%\5��Uĭ��\������y���CmŸH�����;�ǘ�N�>Af^~�3� �Oα<=���v0q�ll��u��/�7F�����ї\����2��}8��T��Q����^�Y�m$Q�is�C��'m������7��G ��$��������Sr�Hn
���}�|�H�eR�?<��C������ʡ9<��q4����Ѥ��C��s��r{g�pXX/�U_	���,I�j�u��f��[���2�D<��;@t�[/�y�DO��<� ��p�#�h�e���>B��������;r#6��ck��Ɉ0a\�z!x8{�MUG] ����mfv�«�*6i�mә^���Sh�玐�
�� حR��`���L����6��W��v�{�~	�B1���y�bPo�j=��Ssa4��Hb��s��6�>����(�o��I�ƊFE�#%w�!R�\ʕ	J��y�q�$P׸�7�cc�eۉ��p���K���5N�dA_�o��ţ~���Dr� ��֜Y��'�i��%���d>��m��sY��5{>����:gU�;�ŋ���b)��|�������CS4�c'�?ru���e������>65�0���an�!����:5��'��/O����{԰�/���ׄ���8�q���p�V��b}������O���(�~�S��;��o��?4ۿ����O���(�f�S��;�m`�j�G�X�����Ql�O������7������6�j�G����?4ۿ���O���(����f�w�?�C��;�m����l��b��h�G�b㟚��Ql�Z�����6`j�G����?4ۿ��������Ql������(���S��;�m0/j�G����Ql���S��;�m���l��b��h�G���f�w��^��l��b���Ql������(����f�w� 3�����6�ʟ���Ql�H�f�w�?�C��;�mЗ?5ۿ��������Ql���S��;�m�1��l��b�?5ۿ��������Ql������(��n�S��;�m���l��b������Ql�����������l��b���Ql�������6�j�G���f��U�m?��b0�J��_��b�����Wl���ձ����Uc����+T��wbΆ�t���A���ʷ^-Q���07"�VY��_�cS�����TF��ԼgE�w+��- H���~�%�o����Ə.'=�:r�h;{=g�n�/�Z�5��@_|���j��'�V^}7�j�1�UaQ�+#L�>7�X�I��6�f��qy���{���)�߈X��3QR#̦˺�~��ϟ�^Y<{M�a54n��֒>���,�Fdg��� ��9����d6���� ���<_�{�`큠��R�Eb�x��v����Vg~�n�Eq��d�)a蘨C��h��*TmO�quZrd戵��gu���1�J��Wu��pBz$U:rIn��D���x>���7e��6�������m�r�� ^*{��S�fr6��NGKh���4��o�{j'�?�����<y�Oy���S�G<{�,� 5����0@�{G
����a+/Z<�E��2��λN�Y ��V�$�h�F.g+�}A�2��XT�.�=L �a7��n�����a�Xz�U��;�E�3}�s%y����\GL��"2�`�Vɤ�q鯩�� ��=��")�!32���p��&��`���9(���Nu;�t&y�:b�Q�́���d�뾌�z���#˃�;ϖ�hˌ�[��Ml����d�������{=�.���؜����k���#)�qs:Ut^� &\
�П���M#p���w����?���[Ń 8��'�mw�Yc�%���(x�1��_۾�f����k=�̂���sp��H�[Q~
��%�lc>���ˉ��u3�o�䧍����]�T�a��{'�j�v8�k���<DQ����D���&kx�)]�_��|���*�*Y����X�BN��tX�t9�sz�!Ti_���'��]H�U~�Ĝ�����4e+?���U�|H�׳i5����/I�%h~Dg��.?֍�pB�i,�晏��1`Q�s'�{3���vi��ğ,S�3qU_��O�>N/�B����/��g����{��n\|O�JO��F'�:�c~#Z���K��3z9:��W�Y�E�b'"������ւ�~���%+�]�B"n�WѼ��_Vu��^Vx�G���EIwȳ&В��ZZ!����ͫ�Il�fK-C�����һ��[��IE�M��H���N��<ݭ�����0����- �N�^<�B e��So���_Akp��}�.��?�p�m���]Y�iB�,�z���Nq7�*����\��e5a@���������G9 cH4��Ln����'����Q*C\V��.VV{#� ?������הp�8�gk{�%��Eƻ���)r	l�1��͢�B���v*ӻ��}�j&�&��/�& ?�[�<�%�Ԯu6�r�4�=�]Y<��:&�hs�}�o��^7��@x봟h-%�F'=�81��I��k��T�7�/ګ:_<��8��<���	�w K��fr���ɽ��W�C��c�R�T��Ꞧ��`�q f805�JG~���a<��!��^�aP=����Җ�:+����wCd��yI(�T����S�iB&7�����R�O��ߐw�αp�g�'�ꇀ�ɺm���"vY����}��%�3,-�,K=�����X�?�76w�i������&��|ڱN�����n|�Os�MT�P���?�C�=���D�@:�#(c��V���CQ���@��[�T�zO���5S�r(kH��^0���bn-E�x��ԯ��{����
cJZ>�|�������
kHY8�;:�oA���Y� ��ŗ5bh6?嵮׊W�������s�$v�w%�: J�b��+�+	]EI%aJ��5�nQ�ԙ�XH����R:�lJ�j�X����S]�EnǼ���zM	VQ�H%r�ݲ}۫�O}�]��N���j�A�ۭP$(wc����%ޣ)��a�����D�;<X�.d�&�8U��t"'������7$X���~���k1�:�;�S���!�:C���j�eo�CD���0oC�yܒ�q}g ����9w����l,��f���T�о�BNQ��"7�i��}`��������?�5��	ڵ�m`�
�-Q�t�[��.�=�KRz�q���Tކ���w�߹��T�{~݂@�d���qȂ�6�`5��YH���l���$�d��z^�lCB�`oF�� �g����
 ���&��I:�_�LjoEN�����M��t0snϣ�g���J���5������-Iܥ������D�D=A�F(^�����Nf�PT�����F ��< ��2�a�b�����>�g�X�[���ͷs+��<�~���r�wĴ��%����!/�}�d�%MU�.���^2Uy��!��_����5E���B��ߵ&�υj�j����\�贓ep���)$Jt+�{�jh��*`/p曹UG�T0����� &'�Zw��}
�<>����K�Kb�,/�Y<�r���D�cլ���.��cd�a޵�K)�ԯ;��G̝co�Rf����*�V�͹�`��^������Bst7 ��h9:��c�&�M�*��%b�'ܔGKʏ@)Pb���&���i*|Mߪ���<.	�pd�I)Z�_<,n�ὗ��~Ϥ<�K )sAt/����lM�#�,�n��$>S�(/1��t��W9�gȗ������~�oh^�kyJ���hW���t�W��o'�]u��C�f6np�H/<�N������xu�'�njP|�#���p�mU�OC!T�g�W��)�}b!ˬ<w��a�����t�Y��/�/�b�Uh�8�?���7��d>��;��o�
������<S�7	�ϐ�F��j�3�klqg�w[�k�?O-��:�[����i�x`���?j���'��QF�3�;�_ůS�DK��3�K��_�~�����r�G��f���:5���?������r��hU�
�����?ώ.��@/�?x>�����˱����yf#��_�6�?��Tk�<��+����ɹ�R�q�����N�n�T�}��]�8��E�65���붓���C��O/- �1~��6`��MT���k�����݀��Jw�M>�Nρ�|Xx0�-�O��7�x�;��N�����JD�;�Cz�e4E_s:d9�s$�d
]�DU�o���la�班����kϡ����2��E����2�Qx�����9Ivkg�Ob0p9�I�@A��쬬��ξ���FN>���=f��YC=����P�Q�Lj��߯pn>v���� �I����zQ90M����C�*��|���:@>���a�BO�KH�� [����9r���M&B�R [�^⎕
N.�:���{�t����K.YC��F�����?����t�dN��+v;'^|�zY,�(F�WO<�GS̀�in��4����� �:��:=Seӊ������Wzoޖ>�`����t�h���S��ϝV���nL^�F�-���(�y��0�ς?%)Ҝ���ʯ�n;��ǻ�o�Ş�����4��[��Umy:��=\������F���pa`��v���
�,��[z=������{V\[hUn �GV� ����c�^��q�_��W#-0e뚜z��������7�7B���}�^	_-����N:G%k"n�Pv._wd:߽�v����}��8�옉j�u�E)ս�8!Agy�T/7L� {V;t��.���s����40�Ā�eA?�����f^q,F������Ec��?R�Ы**��_����L=u+�O��4l��R2����ziV�����3|��&�}$��Ҝ��*�b;�w3�=~BPO���r
��kg��L϶�>~�(�*�����
q�/)ik�F�֫k�~kޱg�YX � N�u�����%!*ݍ5��]�Um{!�7�k��>Wr�#�J<<I���;6���6(�S_�
���)�����J��/8�f��צ
��yc�a�=(��n������Mѡ���f�fx���e��2`��:WT%��gs��~���!�d(�����i��s����K�%K���$�����cQ�(5�3�$�e<��7\��*FMs[
ђ�t�:	��̌z�s�kD6޾ɡ�N��|0~u��Hȥ���%*����]�� ��Rs~2\�թ��o�&92���T`v�UA��W���&%Px"����O��ƃ~�m�<t����5X��R�"�a�jo'��|�7��o�ڞ�'rN_�e!I|��P�ʈ����%�W�����ηk����R�����7��N,�J@�j��H��l� R4u�;�rs�W=���`ŋڣ��ZP��'���S�2p�~�-jX�b�p$E�E��r�d�H�2C�����~�����`�;�[s:B |�
Niru!@��Y)7�l��著;������f�m�w�<��])��2����y���9_GR�7yR�������-(l�"��$���C���a{��ϲ\%v�d	Xݹ~!��e�B����.���D�$�t�]?�);���L5':?K�:��-Y�/�T��Q��Id�>E�2���I���������iA�&J橷17���`��&�y����
�9.	6�`QH~[>zo!���	�ڃ)��PH޷�7��'�[/���Ͳ��ë��<�v�h�8r�kF���Â���RJ�W)4�5K������� *�<��=���I��R���(F�H\�(Q���E$[���F���wG�\7��Js|R.�\؛v������!���v���i�o�F�T��a\��/��:g�/�U��{��#Kݟ��+� ����y������
�GaT�rJ ��1F"�w������&���ղĭ�������:�� �ԋ�@�?ܪ��o����,��.����@����O�h�ؒ���hTag��Kr�������b��
��f� ����_h��S|e�������T��X�����_�����D�?�z�k�F%원��t����ﻗ!T_���;��_З�׉J���10_ؿ�(B�[%@���L}k��#��/'�'��GO����M��ك������#����Vъ��a�������y>��� �Ƹ}s��9c�~���Xd"���A�o������!�v�԰�]�o+�7W��*�k�فchy�?��ע����O��3v���\�������?�Xz>�ŋ/x� ���	�1:\��v�8]1<eu3���|���lB�S���	��m����FC�x@���:dg�P6�.��Y�V��������r~0�-���>��~*�+R8������,���E�??�B݊�N����&��6:Rҹ_���#{YjFM��=hȡ:f�����7��3���
>kEK}����ܿ���Û��f}VP�t͘�O{i�`�X�|������,�z����no�~�H�ƚ��{B(@�
S����WЋ��ڨ>��HoƎ�o�)�4�&��xFNi�������mRu��5�����R��R4<���q#�tzZs�z�#���h�ǧQ-�sJ�sk�tl������#C�F��wk���U�+ػ�D5z;�@���~����U�Éb�������Ӆcaw[���bi� �I���7���.�2T^�:��E�ٳXk�W��/$��[>�#�����߲���!0�����0�/���	�^���=Y��_���!`�<����
!�y�������[�[�v��IK"ͭ*~Ua��X[č�Q�q�����W5��/a����
D�K��-Y���?��׾�dv	�f�G��~QG�%�E����*��N��oӫ�z��0��*5~]�@��g����A�6G��xL����ϸ}���~���������vSk������/>�H��U���S�ei�*-��aG2i��?��m`帙�8����0���,i��9�x�䦜�i��gB��M���v�n���NvI�����9��O��}��s?&b3���t#b�Ñ5��d��l@�ݸ$сM�6�ڱ�Jv@r��=����N@c���ӽ�^/�_a>�>Q[���\�����Q�l1����w��kᇨ��%�<��Y��<�k�ρ�_&���jBu�S7��&���]�yc���I���b4gx�|��e�Dqe�����������~����E�Q���o ����O��#�汜���>a���R7t�4����C8-z]���2l\br�ۄ>`�a�m��I��`n=��(��!*��/��ΕV J8>�~�9!��tQ������/-ȣ�n���Z�k1뀹L��V�Zܿ�^b`	@{f����pN���݁�J��;�;�YM�"�6lÆ���.[ɫ�*��7��ui�1�r����R}?�O�D}{)O��O��^��f���Xu�W#J���������b�zJx��g���-Z�5 �)e�I��-�`���՞e&��(��G�i	&|8���B�9A�ɶ��u� �*G]/�Kmv$g�5�p!a����3�	�BK���򡘧4�~�tb���Ǭ�7_��$ ��c��Tc��B�N��kz�.�f�qT/K��ߜV	=�k�t�U+��AF	jQz͹C���0n�T�d/��X[�����ι�PM�� ��rI���ɴ��0�I��3�Ӻ��\���V����O����:�>ߤ �nz�/�qq�,e��S�� 	��8un���b阃��c���'��`u��|�����gk`۵���ɧ?:�d�?�Kl�3�]C�dg֛�.�'�����B�X�pL� &��C�]>�������41	A_�U���,���M���v�����D2#��c�T��yGA�0�c��p-`^D��z�RQ�T~DMt�V���� ��<�D
��;�IjUD�?^=$���Y'�:=���P'�ƺֽ�᭚Cx-5rF�Yq<�p���am8��k����Ӫ�:@������Zɭsy���A��h����|��{�dyv�&$�hMo~v3I�\7���b7�ʙ�7��BM��{R�RjZ��42/�i�zѹ�e]L�ț�a�1��7��9�31~ji:����`2�bTr�`2�.	j�����d�[�c $��;�9��g��������������K@��N�������������Ɨ���W_�U��Wq����L�n�`���I�����zMv���^1�׫������wο^{Z�^�_����*}_���o�_9�o&��A@D� ���?��}�`���o�u�����+�"$�?b�e�Db���s5%�kz��>���g�`��ɯ���I��l6���U����֕ʀ]�Y����_��G��)�͓��������/~��Lv��� B��ɂ��#�����gn\�����q\1���^ߙ������Ϳ�˟��i"Z�]�Ř:�w{��'���\������_f����ټ�}��q�o��ڇi�;/����?v����_�����4���o����}����G��F��������k��q��`v���P#5^�Il־O�ݥY�P1�_���k}�R�
��"��MͿ*]UE�V��%�z ���<	��#�Wl��ļ�I����K�zQ(�6e}�he��j�&�_�baȀ���l�2�]Rܺ���pg��Qy�~��I��ڻ�yM��(�n�gO� '̶�Ol/�W��S���&w3�YБI�*FԨ�I`�]=�xA��]��4��Ԧ��g�LY]j/+6��*��P	����Ͱ����h�L��s���2+�'o !1�ht.���|f��L�)y�Kz{amdi���+)xq��-�^>=X�a�!�Z��\T$��J�Qe�,xQu�kh����0^��rڠwɸ+�V��b�s���SY+��:`�d�Ґ�=u�C��+m�9��ٗ*7	�4�>�c��|����Bf�q�Km�25F{Ї�}�s�>�d����@]�ƿF���u�\��u�oO8f����u�q`)�Gp(���qj�ifr+Ey�N�2�<[Ӱ�F�~"��H�>V��=3[��4���M���I$���зr����>����6��-�U3k�'pYpߩp� �}G\5!v�;ģ�����i��Nl��z��񇴊���Vӭ?���$�O萮�*o�RF!�i�[�D$�7�*��a_ v	��fx���緷$/Y��h�
!$�㏢8�²��A_�V�3~�H�(���#b�q딚���""��~� P�BB<1��!q�
n�|x�$�y�W�+|}^��:y/)�S?��חQ^o��ߟ�XC�a<}.w@����vz0=�%s�vߥ�0���ni�29�Bz��dAC�U�rq(��k��\�Y5R�4!3rw*���UP�Eb-�����8�'�IEzteY�e��ρfj�텂���{��`+��y)��ڜ͹��% 3!M��C/Ewt�E�
�?p!��i��ZM7���-2�cn|�Q���{�O"AD��G��k�ބ��͛�o`�I���v������UD��U߲�B3�,�08�3ғ5�3sk���#,p��&8����$^S���[������D��,�՘��D�C�!>�������q�V�lA'<�xM}yd�/ �*_� �g�������+qz��=|綝�^γ��Q�Q��z#��]kA�$����l���������$�����Wș�>[����>p���PyuX�CUV��U����Z��ݑ����(*�}�p���eW6R�ى���J~ṕ}�X�G>��������<��{���f�-�+���X����~�����,�7�+]���J('�ݔ]��֚��Cb�>��R%�_�jj�g�$�	��q�q�.M�ܓH�_�&?]QHw
YS^�������?�����G4�'����!���~��.t2n0�&��3kB�k�>�mT�����i'+�[n��-�K���s�� )ѪH7H���z�PX����w��-n���\
I����{��t1�ҹ���������✵�$�ә��Y��K���0.�
ۀOst'&z��|p�-�8SL�*����CP`o��/�i~÷גSZ!hs͈�a2 f�9<��m&�s��ʙ
/.=�Y���@�>vh�Z��SY:a������F��z��3�f`�6�'���� s\~��-�E�l@}�f,�R�-�"����gb^T��nĭb�y}���C�CX�W^.�		8m�/~b?��?��� �n�>��ԜQLAOD�C��Q�I����^�"C���(B�ժ�}~��5vik�к%J�4+���JwN����~��i�x�GϢ����!�Ї�Lul���dn�ֈ�2��ǧғ�g�~�Wcio��o�`�!D5���C�t�z�,W�10�bO��xS_i����wJ��o����Oa{	�pSޮ��Z�1?�1�JL�V�M������?�J�}P�MH��\;�+h9v���Ҧ�>ߘ}�����sl4I�G�n�jےt&4L��������|A�n1�'��c��#/G���>F;o*�#L'4�}��y�[�����kV�����Ԛ<�$Ih���jh�&Q�7�S�d��[(����c^��M��\O]���Y��u�&��}���1!��4o����i�sr�%L�bm�T�^D��v�غ`U�!N�<�{��#�O�o;ެ>�1	��
�͢�Z�ᢊ� F��αQ.�����c�9���Ǣ�?Z1����C ܫ�*����|�.y��!n���һSc���U�0h������^�٬c�\qG)��l@��2�)e���}�~
Zbw*1I�w�Q�'rBoF���� !\oʷ���H=���(7yUi���t�+�#T�����^L�r�����n���C|-I������e�c��l�q�E��9i{1����O-dT�w+Ly��I
�d��!���6*R����R��e]x�xvY����r���Y��WK��m�6�禶�ɸ�}����H=�$�@n� �&C�]�Tӈ77e��bb�qo�D�|V��P���ޛ듔��X+���򝆈��+��֜V�at�h?��P���n��g�z��YM����#�ҳ L�p��$��b��D� ?�g5CY6�L|�1H�@)� $�Gs��%2�	?��D��PɎ�7��p�z�ta�-�A����	Bv���8�Z�4v\��MR���`��!a���H�Vw�2�7��܅�Ƒ�����5�������6��9U�"�I8��n����Z��%�����ܔ�����1)>���ꨟ�� ��hkζXϠ��om���؊�=UaEY�g�L+��jaMq�cA#o1U%�q/�Ox?��V�L�"�k�K�����u/�1�i�
�4���/���}��N�Q)D�y�-\`����tE�����ٖ�PB�+�G�����G��O������Bfd��rV��dJ��S2J����s "�I�DD��<�L�巧�U����+���N;�tx�	�K���cǥ���|؏�|���0��b�hgW"2�F܅�\�%=��5sz��=�y���.ai.�#Z;�+@��թT;J��˵B�弨���9�U�l
��+xj[h���\ʊ$e�XD~4�o��G�#f�[�����#�pKW^ ��l�D(�%#TU�K.�ϋ6�֪c�g#�
P0/��炏XR�c��&�y��'B�k6LT ��#s��G���ȷ_G�6�����o��o�y��VZ�U��gfںQ;�&�?����>0��W��i�2f���۱�ߓ�ü�]?�����bF���|�4
���>���*U�.�T<�ZV,~��������ԗ�u2���b���g�[����m�@�e����V,���?�.����ޖM|�"1���%�O���Q�,:�{����c ����W7p�b�~��`���F!�x<Tng,,e���c�ھ��3D���Gb;�R��>%���i{��� �M"Zdt�� 1��	��#�D�ĕ��fP�46r�g�~>������< F�)} �^N�rZ@{�����h�������/��J��:r��Y�h�ʃ��x���� �|����b�'����6�k���`.���b�u.�E�k��
b*
,F�U���b=��\DdDfd���[�7�IС5�Z�����7<�z�I���I2�5P<��[���n��y�9g�h�a �u�&i��t�4]UK��f��޲\Wp���:맣�^���W���-��"������~�AS���H�J3�8�1���׬2�y���^��G��/�������]�6l����.��p�b��+`� ���+��P
o�]��">��k���E�
ƿ�ZK����2�,����r��z��9�������}��������� K���}�A�%1��rY�9A�dP>?�uqa��IZ}�v|}Q��|3�--�'�48(Kb�E~ol��b͌v�ʓc�mNa��*c��}���ޅc���*Ʋ�����"���zH��onk	���"b �Tg�D \�����LC��;�"���q=�
?=�D~�����,��$���1�����S�3?<l��G_vj5�&�dE-�"�d�# ���0ɬ�V�gE�#5 `tBV!����C)�}�_�/��G3MqR�U$I���Ƀm��ӗ}C�6^��r�GW/Q�Z^�z�.$7����M�cj��
�m�3P����"�}��'��O�jo�v�T����Q�g`o�J�'��'�n!K���ט����
i;�k,�o��;ex���y����q��"��S��s~2�2�<`�p�,u�]���^�_���L��!,���<&]˅���U��n������&�a��α̭�x���?���!��Y�&���vR'���OY��A���қڷ�ُ��J�8U6h�P�F&L�݂>�p6�V1&��6�ʞ�T��,i�!A�L�Zƻڮ������{��
[3��LdnI(�ZP���":���6��=�:�
$��,�����������Ac�?��v�Ԋ ��C����a|����gje8j� ���3%�9�s�c"�|YJ�bG���z��=RW�p�rn<�-��/˒f��栱v����=Kf���V>�"eRs/��K)a�A˔ |��M�早��K����(�ϟ���S������k��^hB4�{�ȳ�H6����� ���Xf[��`8Ԙ-zdb���it���ȍ*�im�W�����$}�}s�����H�Y��*H;���_��~�@�9���6y��m�㿉��[NdD�*S*���z�vh4;�B�D0"���#���'B����?'�E�&�0�s���W��K��+�:u����?Q��}5sꮇ��~��Y�J�R��a�]5�^�8x�F��"��=��Ͻ�?q�]c��sB�3���w��9cr��>ҵ?�[�{?����٘�Dv����e�?'A�^3�?���K�ny�c���ԛ�O\ٟ����߿Eu���3To�����|�z%�+>�ϟ}���;���m,�x�����˸˿}R�k-���=���m��+ȼ�ȋ~��?י5�;�gg��_g{͗8�ߏ����� �J��,��û��9��}$n�z�F�yʞ��سW�Hh�w����=��Y�_�^�2_��z���?�p=�������m���?R����"{?�T=�0��p~"p��?^�9��)�Ϭ�����G���?������!K�����'��hG�� I�0�!tȯ[d�D.RE΋5�W�]J��lY��eD1��1A�ޯ�]��P`����b��ᾃ<}��w��z�Ea&C�?a�6�*jj�ͣ��hb�><o��
CsN�)$���t�B(o2�z<��gf��5�U��O��t��h��ҝ+�Dt$bmCM !_�=h����;̱-�����*�EL���Ҧ�*vJ nQ%�%y�k��7z�G�*<�9C^�l�O�M�S��f��E���c��X%0,}pX�+��)#����n��-}���#Lˬ� :� ��
���i@�ç�^a�V��^sx���MtYL�/�(fA�\�s�{e�1;.�)b���������/Ɛ���di�1�ň߰h�S���q^S*(K��eo��뒿&�p�A�����*��%�4���j��p�Kr�����49
�ч��p���*�N�'p�H�_?��Y������v��Sv��|�&��[�l�{�R�*��O���
/�����z|�~Z'���KQK`�7�e�؝�h���|o5݃�K�-���H���H�íL�:��P捞���ǔ�����-"��2M�ܨ,��(r��RM��ʖ�"�V�P�9~�\��Ë�qP�E�Z{@ȷ�괜[+ >j";5�y���@���A1�����q�`<�M/	�5d��1�e�y�%�J�ʐZ����UJ����a�:u7 ��.S6S�������>����v�]e*Ϯ���.���ˡ�����߿>\�T��y?0����S6������٨�W$V�~�ة0|��q�opX�6?`~l;�l+KR](�	�bj�M����U��[8Ԇ����{�pb�"L%�K�PC�r~�\V�8tc/�V��ǖl��5^�G�H�AL�+�T�3[�՘��}�j����x�m��-����,/�D�
�
�w�(�0[x)=�:�]����#`�X�/�}d� ����<��"�ןk}�m�s�-Csq�Χ�K��O��js����.�h����˼G8�I�wA�����ԓ퍠52�=�#�el�^A	��cDp�[�`X[��zc�E�tn&���&!a~�Fe{t"�i�\�C�cBɒ��e��K>��O�tH�B��-0����5m�z{���;g�>�
my�+*?�f���k�0!��->|�����H.A^V�v����3�K@ҍ��(�U��V;�WE��z��-�S�f 3В������q ��ȸ�S
�:�٬�u7�X��K5�Z�gZ��9Q��,��ay���z�ԢOI��ǃ�8 �N�˃�	�A�l_)��k5b䋢�~Љ����)����=JR*I���5A2�F�!�x�'��i���j�5բPh�9���w�C<+����Q�!d}�J�w㔴�
�{�3��áo���條7�*(��T�2�����ۙ�����z>����O�˱���2����{�@�+�K^R�i�QJzqm��b���$�Q��6k :j����j�����R��l��=|q%R$��p�Ꝕ��%ֱQ˪�xW��K��P���w���	���*�U+
r�$�!�?EW�717Ǐ,?�����hox�"oE��.�N��J�(d��JW�ěIZ����޵�о�Ze�߿`��>t�Tf�fW�6����u6Nv���#��`lq�µ�Rn�|C#ĢL������c��������'��ZS���c,�]��r;Pl�� �������G��=��Ƴ�G�_�i�t��:yכּ.Y�b�	b�T2�UVȞ��9J�j��d��礐�v��Q\_7�Ca��qmy:o/�KO�ŭ�0���g�{�y�x�U�0�q�>x7�GPQ|�cca�?�:/�����EU������\FJd�~��]���j.��v�X������g{r[,���s�|^4��S��=�1/��1��0�9̎��i��d0U\5����8����V����< tuJćC�ے�ǌ�(��_>����E�� m}����0n�Ne/Nw��vr�-Sq����$����l�~fDG:kb�{y�a+�0M� L����Gv#���r ���K�`{��(
G9�{��ܛ, ��l���M�Y�=�1E�0ᑷƠ.�A_�ĵ��s0�"�"~�o=�A0[�,�sH;�H���]��j�����ֶ��oT ��|R���>7r� �����m@c�@��H�
�����9��+��/�:�:�J�Q�'L�5�������2����k�א�Y5�2��Ψ��+�KX�x?����R���Z��n�n����7Ɵ��,@o?���f8S*�*�By�#u���� �X���5��G6�r2ϥm1�Y!�Jm�M����UIğ�Չ��Gk��fq!����#y4z�a�P��Js���T}k��x�K�w�����ch�b��� ;s��>fS�ji$-ʘ��r�ԗ�U��W�I945*����ʱ�È=��{��*71x�S����טjE-��E������9�X9��<��M:�3ݳaj"(��K�n��rJ�f�Ͳl�Z�����P*�͎�QF�N��~�iRͬ� �<��=�^��[�f��uj�Fh���^�������Z��
�u�'����'��Ż̦�5���}�Tk�7*>�k���ʹ�_Y��]��a�A-�P���@���$�ʵT�<�k�I��1�Yʅ�@�g�b҈iy�X�.L�H9�h3�W_��a�!"q�:��VB���݈qet+��.궕s��KXX����UO)�
�}h��x��.�E7�XH��v��m�v����C�h�/����+$������ Gz�0���|�a]���˓}���j�DJ�a¢�w��;ͯdV�"��+����#u��8�cG/�����е�t:q�$��v�T��#nY�� ���j�������r��6����MŖ+����ٲ��M�(��-��sas�m%6���b����b�-g\�,u-���_��errQ�_�Y�^صsT�"��W;�l��Ϗ�fGX0뢝���8])�T�n�p$)uHAԦ2��*�D��+���I�	��y֤��G@��% 9j=I���;x�$=~,�N���vKF.��Jtnڗ��l
rA��߿�O�C�e��"ab_{�e��p�-��*�r;&wO��Z�c!XO߹��k���3���F��m@:����`�	D��$u���e+��l�=vE�6�m��{2�qs@��Ad>J�<�/�ϊ~��� ]L���Z��h�F��#�e<SS��}���O�l%yJ�����[�ƻ=݁]�ڭ�峭r�Ƿ����(�Y.�S]�Q3P���,�X�ܩ�U��4�>��L��i�3~�G����R�U����Ӯ��'F	��U wB��� �_�����5��p_C(Ӎ�^n��t�kC�g�fQ6֏~|#&X�HB�/j��iH6=;dE{�u3���^'d�+@�*��m(�D����xdW���L=Eá|R m��5%��(yC�YK��f5�<�����4 u	��{���a��9�?�*x�I;�KX�J�g����jJQ��x����Z
���mTN�
�|ހ���9c�U;�6ׇ~��~Y����r����<��_%�VEA9�[3������ۻg2$�TG�#�&/���;��Ѓv�^��.����-ׂ(zD6ԩ<((Y0#aOaʁMY6`�?����)��:��%�$L�W��x@*�����P� �YE!;���Ʒ$t�6��8��Κ��~�!N�g��{��x�Y���|�yxs1�c�q������+�v���nt�TS��p`4Ty<..�$S�W���c�$��5u�G��"~���KU���%
�����t8"����q|�(h�0'�Y��˻A=������FrǦ�v�%i��w 9~
�9Kr�8�&�3e{=1�/�cw�h�o�b�\}{1�3��Gd�M@�F����m1!zF' P�0���@#���{J�د]S+x��&S��_U8��0�+�/	�Һ���uBn���h�m�.�lϺu��#oF!�3��vӷ@%]F'}ʨ/���G�_��.����p?�H	��b��N���%�,Kk�J�@�$ܴ�J`3�2a!���G����0�
�l��Po���ˮ��{K�U�8����>��/����b��d��I��y��B1
 ��	Kr ��M��<I�=�<�^��ߔ��rkW�%�7���Ip�$�̱�y��%:��J�#�c��-�������d�#�/35��%Tb�Rv��h�K}��`0C�=VJ0'�-,-Zg.�)p����
2�+�Tj\f�����Jq�}#{���&�5N�Y�8��P���q�qVy��u	��AuȞ�U<��r�êr�H�~I鈐��߿4�2z�ݳ�8= ���wv��1f���J:�C˳�᧤��s0OY���f�63Խ��l�*x[��H��E���fYDP�w�\�`|�hIk��[�	>	����8��x��f���ȿ?Տ'�+�R��1tF_�(����q�qK�Hz����]��IG�y�8����<�'<�2��:r���^��nM�7(z����G�Pз�I�q�	��������"&�qΙE[���f�^��	���2>��D��U�7��q����o,G%JvojJ�%�(��|��?��򙈞�HiK?|���6��s
��-u�~	ȃoVC����#����ab"I��@cF4���
e���5V��F9Ր;|����ι}j���5���
�2���/@B��~��*L��y|����a-ܷ1���S�՟�թܵo���b��TRޜ~)�Ზ?
_+ �?�����f�Ph�xǁw����2R��z�`�y6�"u$D�>�ȺG�m�
[�'b𐸾���R�w�
_|U|iZ�2)���M$u=+��O���qO�H�NC���MD�&_�Sd�W�l'f��NJw��(�A�'W"�I���tW���1�Z�^~Ώ��k�����"I!q��_$�Y���"�Ճ��8���?~�hoX�9�Lzҧ�<��_j����D���Z���ȣs�od	��/���[��2��Ǔ�b��bL������,�U�,�n/�^Da�|{�ey��vֹ����U��dk0���I���Ygי%`�׃��^#�7g�m��̸� ��a��v�b�`�^Ŋ������+BJM#9�9��a��F0���~j��$%L`<�U��3�\v�!4Oȫ�$�n��l��`�	t/��~~i�����ְX���^�*��� R�v�ޗ��	�B�8�0Oc����|tb��3��h6�m�ȬC���Y�h��+���:�S�^߽�p�w��{�^�c��jMfÊ���,O�Q��\ ����V}�NSX�SJ���E����rl�[��'9����iP"�'���4�g+6����1f)Z�3Ik4�+����Y�9��97^��J��r̃�[�]F.�-��J)n����N��*68�KP��!A��F�;���~r
}�9�W=���=(i_*��g�4j����|M�`����c�g[G��t�ˬq:�A�<�")@���fT����bn��l~��{��@��̿�g��E���+�i�Î�����*4���ݯ�l]_�(W/�f
�v�.*�x��k!�F6,m���F�+}؄�DaJd��2�y~�T����_�HAl�?:�/��+`�,}�nӬ�_L�B�N��kص%��������X7O�ibrDp�+�=�YI��0�����y�Hw�+�~)��Ge=�@�H�S�ZIA��q�#(��m�P�>S$Yrl�{����.����C2sQ<v\|�\W��`�[���[*k�J���h�-�)�x�� ���{��4S� U�NG��p2�"D32����� ����t� <�{�Ի�S�D^�G���
&s��)�˔���� %���ހ�<3�q�%�Z݃>�@���y l;���ƭMV(�p�Dj�:~�!؊��٤�(U�).��7�T�H#9���(�,���̡�Au�#/�q�:S�
N���>+�F@�"�EW��=*�~V*I�����Х0��*�P�	�'
��UQp�Pƈ)��=h�A���
1�ex��kj����t|�f������}��_"��+�ԙy`{��7܊��������(5�%�e넂a�R��0L�j����I��x�i,� ����T߿.�����g�.�ۏh_�i�"L��0��;�Z�Yo"��N�a EE&��������Ut��D�2��Wߣ���S�HP�<�$� TQ��Tz��#����ϊ1�Ai�΂�۵F��j�B��Bo7R���o��ے��&x3�F�{S�n�-�+X���ԍ�{$�?���h�	�.��-�}4`�(���@X��=���hC�)c��������ܓ�ʄ�l1�|�����p�&~�銍�v"�*8~_��ąG槓,m�R ]�}H���..���$��Ra��"�O���<
�$�3�WWB�|Gs+K^J>�~��%+=S��^��������%(�s|(�{��r5�����-&�����id�~hΩS�|�Q��1�
t��v��ȩR{[������q>�op�.�!{VŖ�N� ��)ά���U�lX�Sm�S)�U+��Z��N�G��n�D�јsۃ���NK�r���f������b?n5����j�?�"��3�G���竹�+��%`Tc�4��N�<��]S�Clݮ���u��u�'M�p�ޮ�C�}x�m8���$3e�;Tu~>R="�t�Õ4��@�}}C�"�	xG��={Ē�@��<�p�KI:5m|�Ƭ��C�Y����(j1���i��I�Kd隧7����%S�93"_��b�[�]�jJ��/G�"��[=����W�#:�!�߿�N;?5혵�f�7ue���Sw�1E�eL����`l���@��b���-�G��.v�0���b%l����U��p���:|<�OW�`�_���^ǥOP���+�O�ýB}l+�~��N�9\�i�ʫ�{=�[�4�AMȪ�K������U�=��<���y�)��EdIYUU�F�|�9��!ʃ�������@����$";��}z,�ɔI(�[�o1a�%r�W.V��k���I��{WV~���h~&��F�y��� ͅGj��*-�R�&D[�v���ֆ��Bõ�g���SP�B�|�V��K�'��\���&!ƺ���x;���zO��7�W��n���ݖ�~
3�<�� >�gF�+g�r;![8/�x���8px5�V}��BCa�<aUv�+c����֫�}k�=�ld�����=���/��'�}^P-�IGE��{�%5m��8�&u
���g'
m1;y𮥺����������MD�z��u��2�ܠ������N���d��C�z���:?,Z�ǂ`��Q�������^k��w2�(ټ]�a7`���J�w_�[�{����_��2ɂT�+ޥ�鹁�QB��״ۅ���������uc�: �C��ͤ��?����>�
���q�ޤ�y�8��}[^�s���'�p6^��H�P����E^I\�ё>�� ��X��	vΡ+ʍ���l4�O�(/���Bd�k?e,}���>��>�:�R{ƣƭ4�q./±A���b��p�$=�ɣYb�6`j�o�=<���ŏj��
��{�|�K{R5c��B{'D�i��h�D���}1�� i"��h�J�\�yl#/R,*�r�ҋر9��0������t�pTw�ۀ"�	.�>��F�7H� ̓1���i������YL4$"�(y�zS�y��di��7�^����I��<> �^��>I}�7_s�?��G.��9:=�X*���MZ���s���i����'o�y<�;�4�)Gx(4��p�d�%R��0�2��cZ�֡U��Ą4�{58'�'����v�v�Ko�����|�=�������i*���}*V\��}̱Y/�9	�z��a�N�F��B�y�<��1_7����7C@�`9�a����%V/Zx����B�!�Rm�Ԡ�N���z�lvF��ҏ���V��׾��2��(46� @d�߿q���F��d�^�c<���f��mV#}L�0�]#WH�҈N�0��M>����ש�h���U�H3%<��W���.w`y1 E��2䡤LR���bؑi�*����(#��/���dx����HF���h2zɼJ.`t�Mf��JF�	-{1�G�YW��b�������ޤ�!U�6��ޣ�9ZW�UV�TƾM��M+�߿D��%�׶��[���t��TV9���A ��\˭ϗn���%H�j'��??��/Ex�L����wչ��/������~*P�Q�w�"��	Y(A*3	�0@*�i�Q�������'����O%��[�Pi�|��M��*F�R�e�o���*V���?Yf�+2~��]���y�7Ǜ�οf!<�wP�S	?�_������`����?#��\ȦX�����kp�\�>��Sc�G�E�-�U\�4y��U�D�O�?������[�������Q���៊�E�������S�T�K�@��5�����W���
����ߌ�_s�����E4���o>���l�~���י�kd��i�_���{��á�o���X���z�_��_��ϊu��M*���̡�*
g���U/���:��ײ��&���K�s<�O\SB�&��?�s������?r��&��G����?�s��&�}���������?U��з'@�݀/��{Eߧy|y�u�����e��	+���YYƲW�LcU1�#m�����Ћ;� �z�;_� f�n)�?���۷����}M�q�� �[����L�w<� �p$HZ�nH��@��]P��?�
�?>�V���gڃ����E�a���|A�� �)|G�����K߇����_
��D" �C�L<%��2�z�D�{��
��g�أ[O��w��6�*AD��KD洱�4�pX$dAe�[��IM�WN�C�`�xT�^)m����EV$#q����)�~�B�w��HW�o�ܮ��Xw³��+ �@�.���3�2�&�\��0F8?_���M]_�>��ʠ.�����^��r�d�/�$���V���"��{С����v��m�/9f�w+=/{�u	�	O?5.��V�>�i�����0���)����0��7D�����Ѵ�T���_!�7�<�C(���
~��K3Y�<?ڨ���fuj��R.;Zᐠ0��n�,�ѕ�W�[�q7@I�)��Sg7(�D�Zd�� 5TO��]ea�F�gO�]���3����m��"ϝ�����p��TT���]8Tc����^&V�*4VD�\�0sW�yjY��*Ut�$x�iS�Ǔ�/���S��doiaձ����8�:�*�k����=��" ����D���=>��xE��=@�!58�2�5��9ubW������;fqt^�c*�I��u�k��qz@��a�T�3
3�R}K�l"��of��Q|��3ն�,�<q����&/I�s��~�2��|b4�}�����{MV�@��U���s�/m�E���/���ƺ����*n(ri��s�H��zk�)��{��	�vߌ(k똿r�M��GzP�O���ZN�^j�۶%�ѳ�y�Y�w^�|�j�ڻ�Vm�n�����������6s��Q�6(�ouԷݘ�*�7�N�^4�Hm,���s����2���\6V0���S�|�W��.�Ŷ��5��ۇ�W<�E��hm��z��Y5# z�f��L�e������飍FF����D�e9��rU�th<��s����/�,����������Wλ��\���Ca��p����﨎L�Q%���=^Yʻ��ޯ���Q�߿�u[[��]�Q!�٦u�'Ʌj�p.�ы��,c�Qϴ�v��`X^��xH+�� �� 1��F�!�}�m��_�7�]��r�>.yv���{1,^6�R�/ ��c���̣�)'N��^Q}�2G�8�>�4�̗��ՉGb7.�'sD�}sC/��Ǿ��l!�l�7��}��[�B��ԗ:��b>t�B2߂5�׉����U��r�L���:�&�Ǚ���'�L�tP��j�����ĻgR�ݵ#���
^�xS�W����|,C6*t"����8y�T[��&��~�'�����W>ڻ�t��a7�˳��x�߿p�8$Y�0'=��R��oJ�_FL��K~Q��z��Ky����coGS���꟬���q�P�o���^G"^���pB��s/l�T�Al-8��u��t��{0��%s���H��.?n���B-�0��^��h@ jE+S��Ib(��0����b�$�v��s<�Җ�u4z����%�R��x�:tE�HN^�@=�J[�:��e�KāT�m7az��������P���~��mP�K�#L�Z�=]�Uʽ|!�'c�y6��Gl��������m�AN�Ģ�Ǐžѷ$�[�t�g���ǳE�]��O��;��Fؕ!W���J��OHэ�hs��_{�C�jQ� :w��[�WDP�#~�@&����k^
�ݔL��p��J��c��`*�Pو|����� z�~�b��O�*]��D�ڭN�e>��B@��hUŐiD�mH�sg:�d��)�
�|�����5"s�/o�V!,lP�`�k�h6}oW�'�6m��Nt��ۑ�!��D��*成��+D�'�$|�pM�Ψ�`K6Z��=0^%�t�Χ�Q���Ve(<��DxH������1�߿ȁ%yᛜ�Q�D��za��wq��	d�q��Nr���!��|�[�Y��a������z^H��q��e�Vv�Щ��<�5��28�RW�hW�.d��b@|��bF���tn@��ֹa�!��v���_T������P��u�}6����Q��!y|�JH�?lLo^�i�Y-^!�q^�\��֓8%�.r�R���IE2.n�''��y�w�c1��.�%|�k��kq�W��%B�z����x�:L��E^we��,��C���Aey8ɸ@9G��ݿI�^�i|�f�#G5��p�־=yNߊf�Ij)�QZE��:�?�o}x ?������LK�n����Z���h�������a}�[�LO���%�1��O���247������+�9���@_,+��6K�h]6�Y����e���Y�VU�ɞE�5�6N��3�?��$Y$\O�/�w��]�����7x��֧�!�Lym㟘6+�F�f˫*OH�����)z��޵(�$��f����69�����n����Y���c0mշ��Q��G�BA�!�Cd\�;��!�eP�v����Ƨ]�Z� ���zY���<n~L�(�!���O���^�<]Wa5�r��3.:z���e<�e�J����͈X��;Br"~�͎��;�`0-�u�$�{�v�|�]����b �hW��n`1�p:�;��^�עy��QG�K�X� Ґ�����E���?HY��#��D�{T�qn-0}ǚ6��D�g���<���5Z��Y��,���p��4��r����\9�$��ܦ ���	C-5>p�����hŮ:���C�T��Fq���j�SoW�l;�}���+��/�h��A���=:�����ބ��#$w>����8��:1�7��(]���H!4R��+�@���,�b�5a�bJ��9��$b��#b1K��l��$��o��_?��d���e�h�6��Y7P���r��0���c X�I߄ǝG+D�m�ɕ��p���j$s���'�k�w�_k�G�&����j����Ԡ��A����$��(��"d��Ƈ飬��s:�7u� 9'��_�g�D#���!��ى����ʩ�nK���8>�DWa}�M��=�E��`>���iܻ�����E�^4�����x@ݼ�b	��2�x����S�c|[�r�<�~�}��K�SR�+������Q�:U�uv7n=an^{�J<�yP�v����?\-|��n.�	)��*>U#[�]h`���6�B�h������1��0����U����<Ji�	��o��v��M��e�~;w�O ��˞Q���Yһ
�l����-��q��Țć���%�4l�T��f%<����gi=D����L��I��V�y1Ki����*��ҮA�~���<k}���Ys��Z8p���Yn�+<�3%�:�/kA��g]��N!�T e�w��I�q�!l���} 9Z�!���e�7oj�G{�>P(W?-���ή|IsO��j�J���X�G����k )H���^�8?V&�@�̺�,c���2��zn�͇)���39"��6'�!�k�T{�ul~9$�%^B�g��'z�(�93r�����i�[�;ꄹ�<XH`aݟT\�z�W���
����X~����l�ɠT+���0X���à�?<DM� S�,� CЇ��9^�$�An�QR7yڹ?(�|q�p�#ޟ��mOǓ�J��_��ddq��ϩuӨ�.�;���/����Z*���M�S��D㓊�@�<��?E���>Z5ߚo-��	B=�k{�zz�\�N~l�:o�+��K{aS��_D����`��+�Z���I��X�hv��m�
_QQ|t�]S��E�PQ�8��ą m�\H&|���}O�Ry�{^�.���H�A�eWp�;���=���qY>��U��<L��x!���G�|_����dU��� �u���b,E>$g����9cgʸG�<�3ݬ�1t��7��DD�Rcz�oXC?g�&����Pצ���k��k���-��{7Y���Z3^���"���x�C:���MA�����6v	엺5�����,�\T7N��9>R]�z��g��*j�9ݻ�p�����
��v51!�O��t�l)��ɥ�ǿs����',/��S�BW����p�Æ&��:(�i�X�V?�sL`�f(�f$���uO�HJ�;�X^��p���sHD�1SZ잝��_S(^��)d��^h����&��3_UfZ���!��-�v�F�ꧏ;9Y�f?��ӭYd<L��hY�/���]6�������)����xʼ3Ƿ� �3*��I�:,~�:5V����s ��I[���k�,�m(�r�j���H�w����>_�m�3����٤�S�d�YT��N�V"�u
6�&�"�	�Dƀ�2"�2'���A�RO.C�^�蝟��Nj�nD͌�|�ό�u3K�I��OJ�z�Rj�<���~��N�����g��J��6!8Dm�&�6�X�{ch/8
��M](0�%�M�^�+Q~*~~+��?J���i
�_A��������wL���!LPo~؀�`�P	r썵�|�`�b�D?,y8�;�M�&����Sa9w1���p['���!������Sk����x&ɏ'�?��N��M֕VL�I{�㽿Ѿ����|S�F�90 N��Y��F7��K�['1��IT�xQK�D�]���V��tމ�B��|��Vf��p�0�onR=��ܑ��A{��i��lb���A�e��xq�|]���^������ U�����xfD�C��Cwʋ�>�h��r�oA�6�<���7%�,�a$�d�����}ڕ3�����hh(���$���<�%,Z��|V�mZЯ*����{q`*���
\���tk���T�a	)�Ȟ�5��
o)&[��x-{���҄t_��j�L� l�֜�@��@oC{|@� ��x����;���?wXmo�_�+�s�d�����������O�;=�����9�~x����-���� ]����x����9���I�s�h�ʞsl����J"���?��8�i�?��^��v��O#�^X����8��P�%R�eb�D�%��>�U2Q��9�`�>����37�կ�t(3��
?�����笘����A�W���^��%�%���w�������r��ə�=���S�9]�[���������3��q,��7��k���7��|�	���ߣ0��w��ۿTD������E-�������/j	rM����g����_�l^�����_���3�������O���[-A������࿩$��F���:�h�ʭ�}�Z���WZ�q�pI��²����QV�Ǵ3��6�a�<�72���蟷�}7Up��/�_��;���CQ?���44���U,4}�{N!$:�h��i�7"�+�7. .�X�V�
��tw����<� x۟�3_���o�*�c����-P��ūbƧG^9���'Q�W���tR����%�x��t��=���Z]����^����"L��ѰTo�ą���Z��������R1	4pVf����f���_?5+by�����^;��)i�a�,��QeyYITD@х�]4��c�5�2�G0
���Y�]	��6���Mbz��z?�y��U2*C[�TK���1q4jgŕ5ʟ=����yn.���}�S�[!7�h�1қ}���[
���0Z]�I���p:���XQ������ˆCEx�ya�l%Q*�ex;�g�!Zˤ�&�"s���r~�*a����KJ@��k��1�$"gy_�o������?#�&H�o�Vr��/m��*�Ι�F7C���}}.%&1����#�u�@��J�/#C{m�y�e_��R}"��G�a�VnR���9a��Y\�
�l����T1�BL�x`Y���P:�l�;Nå#�`�j�:g
�*��>��w"�ׁ5T���y͐\�/�~f��Y[q�1K�[@� ������@:\�1j��������S5<��b��\S��á�U	���BQ~9��ouA��lڤ�*4(NM�z�}˴��x4�}���~��m��	���߲BGl��O�G��.v	B惪�:9�sb8�=D29[bk�2^��p��y6��b�{�B��|h~"�ejHo	n�[h?E gM�x�EzG�4�, ��9��2O�>1d��?���W/�� ��?�J����D@��y
�50d2���kd�8�хv�9���� ]U�" � �������_�W⠞��^���Q�K�� R�(�IJ�;P��������{�%D�m�9�A�u
$�1t�>鱦R��+�@f�޸&%X�8� k� ;j+�9*L��)��:�mՐ�2�����u�d^�{��4�w�J�y�����$8�hHB�	��P,��F��o���5���Q���qn"�~ �ϷWI��F�K�M�KQ� ���h�-E��W�4,H� QUQ�ʇ����X�I���a�����./�J���ka7U�{��Xh�� k������4I���*���Q�N��u�5Rɪ�� 92:�(f%Xfl��m�5��N1���w����$]������h0��R@����
+eQ֜�Q�����
Y�PY���j�`����+���Ƈ�D�wl��C_����O揆������ۊZ�䄚�rU����b�6��^��(_3��Cم,�?LxHY�b��i��u�
�C ����Zu�n����G-�*��dh�}�������Z#��兘De�[k�4l ��k�d넹񠤶R�dGQ����6��ǯ5����#滾%p�g�;^�zJ3��҇̀�E�z,��s�4��ؠ��c�O�>�+��3X�~2|����%���s��b��6\������߷�G�r�۞��4�xu������-,�����kE+�i(��t8�t��Ԯ���X�ug���ޔ8<��i0k������/��g��y[�:�sG��hSL�CH� �K8(y˶�:�u	��.eݒO<�\��HAX�ϫ�Q��Th1���	��7{i���gp\�nVo�^Rm�A�����K�v*Kݰ���2dO�k��JӨ{��w��֠:�f��rmh��b;2����?]�����vj^ԝ�$�#$u?����P%���F���(!��p���F����iY�qϺP��߳�+}u�v�1�������vo1����|xcD�>�XM{E�c��?�5?�Lɷ�X��`���A��H&�@鞹v�b���qTn�n���p�R����g:��i�2���<#���i��PPV����$&�J�}�mlrb^�+����v��u(��*S��o�����$��n7`�{5!�
����@����N�D�{�Q7��% ͌;B뗃~����w��ð�
�{c���m]l�V�@^m|>���(�:}Ky�֛�gt�.�2��K�Zh�U����U�>��t�US�j[0�"`�����빊$���q;��sl�r�(�0���b@8��h�z�
�p�R<�HT�K~|fħ/<*#�������Ȉ�]���X`�9-I>�Th3���@t�P|�A?p
�~z���O�	�Z�����|�;�O������>�é�{�5�+�*��M���0/�a��\m}��_��� a����EdKvi�i;F^�*���Ux.qY��`r�pp�	�\� 2��y:�!�=����&�K����$b�㧾I�}������bds-���9BF7��lʎ�o��RUECK�ʇ�������b�ࠫB�6���,�'9���1OFm��8,>-�禔���u�X��<{������;#)��&�'>�������oQq�z��=�%bo�#tXG�^� l`7����飻�p���k��ō h� {�n�r@��}�0=Nl��AVjd`��L�13Y�;{��h��OEa�P���z0s�S��(���O_�SK&�����긓���׼�b�=s{,�߲?z��3K��6��@�S��h~0n �	��&q��q�[`��D�s��>�@<U���4�f�1|�6��c�mQ힉0�L�Yi|�^�?iQ�����ɄU[�|�:�v�\�[��c.D=2$벬1�db�F���1{��e��v�.+ʌ�������.)�����|tю��D�&b�3�Yz�냦��_ȧ�a�#8�l���5�`)&�a�֢9A�+���/�y���WO�����%�!@�A2�I7'(�i�ˢ���dN,�U;�����0o�������ڝ�i���:<=W��OJ���`���K����6?9�ӭS�Z^��+d�wp�q�?>�v��1q��抟�R�1�G�W.ƃT�Ĉ�Z�	�C�@��\��ؽ�mn�c ˕7�M��.��M���|�P�����,N�V���X�"z�Z�i@�)�|	jբ��&�6e^/�cD\�AH�̈��Iv�,!� �	E��a�/�e��.j�v�������һ��>�ѹ�t�� ?,��ޫ�������}!��˼��T|sPhܲ @�D#F�N����u@"E�p�Sb���#���d�jE�`{� Һ0�IR*\a�SRϸJt��61�>�)���*桰�(:�B׀:�
�Tp�{zg#���fe���l(J�f̍�$�M8��Y"�a��������*��N�0�)�. `Y0� ��C�� ��3��v-�t2�Yl����6ɇ�Ŗݴ�@�QO��x}�x�*��������gm�S���Ҿx) ��ȃT�r3�:rQb��<�,�,�nI>(�V��֎��&�ٌ �n���.P���A���`\;3X��E��Op�8��kO}6��kH�����J]ٺq��)�����h�M;q�U�w)|�SPY<�n� ���_g�� �@�xg�a�Կ������IB?�g�� ���b�7{�w�g 9��|܀�#[*�|����' t^�h#z�>vA������!����7��%]������:��C�r���l�b��FB�?����Oz��%�k��|��<�_�� yD_m����2fu�R�ZG?�'MQk���߿p��_�nM����m�:��׺�K�B�%��x��WP���N(��8�3#�sj��
�מa�Pj�K����ʴg��}��Ϋ�F�uS����Z=�c����*�������4,�䧰CGc��z����E��<���j FS7�ZU���v���a��F]�s3�a�̛_�E�u8� ���U}m��Ey�[c��y�t�HC=���ʾ2,|8��.9N���?�4}�>��Y����5�e2�3�Ǯ{\H� L�,A��-�\��J���F����9���7�|k�*rM�^���)!�-��b��m߄�����8�&c���K [V�˽�o՘��2��'���lN&_�Ñ_��E�U����\���_�@��w)��W�$�ͦgM�]م����+�)�Q]aZ���������<�f[NƢ��G
��Q ��i���q=,�@tU�)K�� qTc���i_+��L ���$ >D���Z<��L�#�rDP=����3���\�e����{��05{�|Eŋ^�k5x�����ſ̫�j��J���&�nQ�`�C�Ha��S}���1K��]����%�f���&�q�:���MŁ��ř3��28�����o�K�*|
������a"Z�'>�Ĭ���n���N�B=���� �!���	���fİ
����~���	��]���Ť�����}����s���{�����8���kK��Oa�~�Ku������������(�~J8�NJ�ݶ[3S��f��S
5�3��V�T���T(!�w�U�ڵ�DM�&9HcXaDh��h�Bv� �q=�"*�=�jk�~,f*��ej��*Z��`����.��Ar��/�M���r�UI^�C_GҒ���W�Z�앾�9Ǯ�T�Gc� F�Uq��o�Y��RV���*�nZ���^7��w!v�Dŏ:�S�Y�j٩R���|V�[�f�PKc�f�?C�H�R���u��a�y��ߞ��� H
�un�;x����Gނ�@63"w8Ҡ��tx��i��0@>������/](z����]Z�WV�ӥ��-���Q�����],�����T:(���=z�i���	3������0OR,>��jŤ� YH�E9�2�W��~Vv�O�ovD2�oV��4�#����*<�5�ّ'5�eŎkT�O؞_v��{���E���e�)a�z,��0���7#~����ȷ���y�q"�f��s���L��9cOs��B�ϟ:ڛ��%�ߘ�z���i��~9h%��lo���'��<��xZ}�ܴ��H{�*�+�y q�j�.l� �^.�jF�C��h��K/��!��.�b�K�[l���p�������Ƞ�s���`n'��a8$(v!��|$m�]���&���mB��%��G��j�<�("�L=�3!u_%������j�,��y>(��P�jUǣq�pT{��_,��<B�������M�̇}Ӑ	|������U_c��!��إ�X@��a����%D���9q}�vjM�
����5gH�_��=��E4<�Bizxf�ߨ(����T#�Ze�ݠ�����Yy�����F��SY�g���{�;���
���j����I��U�d�]��G&`�Lq�m6~G�_	�����#��e�?,�[�ʥ�m�����]���㶳G�IA�d�8���2S]��i6ѵ�}=K�\�a���y�T�۠@Ӻ��?"��R�
�ֿ)I}2Ǧ$����^!}���nW�u�?�"�6+��y��8�ho��P�{���v�"sk�k20N�W#/ba���%��5���k�)W�4?�>@���C&���6������YZxu��M�`�Zʃ���J�M>��kܾ5y�L,(pk�g�=!al�E"�&�q	�T�:�hm4�|E߉|_x� ���œҢҨ{�|PdL��jy�q�<�5	�w�0����� ���+��u�{�`���iZ}�];5���؟��tw:�&����N��J��A�����*H!>j}�p�=��W�
��;�RMx���-]�B�S�ed� �.�nN�ٓ��c������/�����>|�L���t)��w�
&=���&�V���U��˫��9�ޯ(��i�5����=ǂ\�%���p�[A�
E�B?%���@�[!�ȱ|oOӦ�u��y�bk�8A^#Rll�)��!.I��Řu�x���1c1I[�¾lě����jm�A`�̖�`��[���h'�@�x�U�x�3����J���n�Y�|u䧦6Oٵy�h�ܚ�Ui�3�:�h����_�m¡�`��%*�����"�`P��5��ܓ���7ɸ��]<���>��[T���I���s�M�o���Yb>�.1n���}M�O���(�5����%+�7V���>d<6���ŵ����k�4P����Y�Q�*G�ɾ�w5�⧍�z�	)�,g$�N�����%V�V w�2N\�v�>��2'�DK�/oz�H�����8L�	BV��*�}�F9g��(�;���%}����I�1ϸ�L�G���p��M���:�$e+h�!�l���*�Tv��-+�?�d�=��ז���伿�&��щe��Wa��6�x�.�2z�4�l��3�m�(�q���oѻ݄_��F��;�
�p�u%���.ύ��̼��%B���O��H�w�G�$�#��r���sL��A1s�&Ļ���B4��S=�l�I����MW=.C��ϴO��wkB�"�E��4��^M��\_��᱙��K+���
����/�X��F�UA�"
ʞ��%��|g_{SHI��T����� �;�=
J�ޗP*�u�u��Tipa���(�����Y1ɏ.2M�1;��iMP5��g�T�b���\e	0��g_>�L���(��2��q!�M] ZNF�s�ܤru�r�9^59+������=W�SB�W���kwX;���� 0�;�P�p��΃A���1΢\����>l�ZǺʏ����6���螮�U��.�o¾�)<�/k�t�H�u�9L-�����L���>������� ��gp�L���)�u���M׼��u�t��Ȱ9�؈��V;3���Z��j����r��r���D�WO�uB7�����&N�ǿbԪe�<3c >I��<�/*_��:��C�!�HmN�(Y\�E�aqzL�q��Z	1�'��Y:j�M$ng	�1�\h�8��a�7�E|/�,WU9ۨ��q�%�����t~�T�i\p�Ph̰��F��1gU>l_��������|����ޫ��z���+`��Oqo�A�f�0�C�)ȿ�����!�@i�ԤW��ܵɨ�98M�W��G~*}l�Ws4�,_�h��N�fsG(_1S\$��Vؘ[���r�oSYk��`���g]�A����b��j����*�-�cU���h$}�l�������_9���X:����ҁd-_x	���R��-o���R$B:0]�:mc���Vz��o��:#}'Q���Gv� 3��f/�n�q&zÊB�^��-�LL����⻂��Z�S�E3y�; ��G��� ;�QT�
:��[,��-B�t�71Mor�wɳ�o�>�	#�����$~z�ڪ����m��D�{�g��hK�ťK��
C��^J��ʰf�!h2ת7����0�f�F�Qb"5|s���}g�sp��Q�]g��}��Ȓ���{(fXթ9��ޣ��cm�N˛�d2�����h��20��9 ?hNkp8̱cf�������:��s"I����1��}�e0���8u�9C6Y��r���
���P"&l?Mǜ�-f[q�Ly��}_*)�"$h�l��2Q��İ�� M�Q� pj
[�0v�x,�"��:����־�F�x�K!�TL�H���7�P�:b:�ޚo\MY���#�J2���R��i��5��t��E�Ma(��Bou�&�ᝏ�>��q_�������?�j��n�^5?��xˀ�'Y�`U�f����(�/\D����༸���|�PÈJ��uW�u��@7U'���9 ����`�	,�s�,g�C��K��f=^���"���Ot�%����O���Y�ڬ�Κ~�%�0]E�(b.6��;�nW贉_ڳ.~=]�z^��(�Aʞ���l�/���ˈ \F~��+$�D@�O,�ŧ� |8�'M�*4`J	E��?2�#R4 �>�m�'��0����)x}����?{��o�'x>��c�.�+s.c�K�FHl����]����� �QȨLߝn}�w�u��AA��굲K�W�g��E*��s���.�G�w}���
�\$��T5N�	NQ��OC9�·�l�dhby�����dr�Pl�z2�O����(�3��g�!H��-�=z&��	)�Uf��l*���>|���ի)͆4k��tV�G��a}��8S��JeI!���Yt��33ߵ�1Xp8�h/_FX���u�W��@j��23Y�R��Z�_�̭z+q20�d�+�k�\��R��V�x�I��^r��0$)f#�n�D=6��颦R�/#�+��x�t�
����1p�mU���txߊ>^��b��j��4�'�8�7Ű\�+���.�c��PX�AB� J{��1ͯb�ף��B�8�� ���``�e�=������M�_r%*/f�#�ِ���7P4<~��[@�D+X#ݏo�yA�����܋4AՉa-IރO��|ʥBE���
]'�'P`:L]%�窵~|#�����I��e��n~�#�S���NAZ����}�D!Y(���"&���B������<pVaM)�1>1x�����n��i�a��ʟ؛��BY��fM3E鋏BN���}j�{�W̘:55�.3��pc� �n�Q�Z��-%�gY_��
|!7d2���f���Z[CbS%�l@�]�q��i1}���A�}^�L�� Hi��S���%��	���`�eH�˴���q�T%p���-Ze������`���s^=�����Ŭ�؁C�&_��G5�V�|Ĳ%�W��1t�!W����������[qwa?��z��mb�s������>
P�4��F���W)����y�G�=&p0�L����{���]Ŧ�xy�����|cՇ����G���gD���1�ҟ�$�~��_V͸"���\� �@9|���v�j��&��  ��h�BYZ�Yd��Jl��A�E�4��4���Ȗ���(�k0G�Y���`�����E	�=���&�R'I=m�
=d=�H�L]Gt�~���vm.��L�R*
�xG�I��#�~�G^̡X��v[��z��[ ��a0�ɘ�$%/�n�%�>>�і�g[an�>����Gvs��8�PP(	Ea���k�������X���2���d�h�d�m#���^�~������?RA� s1����=��g,�d[f:��mNcLL@�� /��EK���LRJv�#c@?SfbF^�#Vc4L��rf/=Lٱ�[6�����S�j
8>��9�V(rR0�y�C�;��E������B��ܳr��i����$�~|�r�|��~�>qK
I��Z�|��h;��v;5�b��^YQ�ه�8Գ.^G��/��nr rv�7QT�@e�h�03�%��6��}�Sv����/����6�����C��_�_/���������ja�aV�/O�A�����8�(��O�.̊6�>���}������/�9���3��\��9_�q��:��3����f|���d|�����dn����O���:�{�ؿTj}��/�[��JM��-�_���yX�z����������9a�������(�}�o*�>��?c��/���i��o��d������Oc��;�����O�T�����_T��k��ʥ���oYe��?U\�?��=|�?����]�I���b,�w�*S*���'��G�����Ez�����]�S#uJ�������6��^������B�{,v[��ރ���zz��?�9���}��Z,�|��~���+�a�����3�;�3�Dzwi�W���:����.^i5���Z�C�p��A���ֆ�i�t�֒;�ȅ ډ�me�ǓYN`Ƕ-[�y�,�� _s��z��u�����è��f
��L36���|eí�8�H�+��{G��b�A�2������~���(�/Ddf��&��?�#��3-�C�"�v\cx<�p"�(!ٺ�<����Z
c9��_l��a���Ъڙ�p�����pmrw��ڟRyq������\!/����]-�9�K��lZR�l�N�4��OcYb�Lɘ�8��P���/�����@{|�7�N��T�^�L�Nv����\�����A~����w^�اq��
�r_�$��y<�� I=X�N�'��0������X���x ZeԐ���-�7�jb@�	)�C��8���_�lo������_�)lk*��7��C�Q�p[)�e�/����0W��KIX��ax�Sڒ�z�Lrq�X������F��W�5����kP���%�y�G2N��	�������=v6�0-������\�X�I7ϱէ�4[�`�߿�pKT�DhrF�Et��p�QF&��'�$n�ޱpE��S�6>|���}7��OD�-��%��Hy���z�+�B�bj9~"���۷(P_u~q>i���Q��=�����rj�ѡb&���e~�y����zZ��Zꬫġ�	HEv�8�:��tis�(;�檉՜�s�<��a�,$�W��nGI"���p�^�����Z8f8N��@[��3��V	��r�9���e)1��U?�v# �F[�̻��ũVuwQ`��_k��'Ы겁Z_{B����WѸ[M:n�ƅ$:X�S)D4_U����u�&���N9.~���y	3/�K��6-�ЛZ׶�P�k�����[�*I���̧��Rw�y8�O��<H� �V�a�@���~��&�Ů��3#s��U�kwD�	�1w>3�ݐ9��^t$?%�O��I"�r�wg
Uʂ=���<S@��F��H��.�Q��O�]�e��!�8������f��tP˙8�z|7K��2؍�{����1�:7��-Gt��0��g&WI�>T/#7G~^$���X�(�� RL����̎�S�W�=d��tD�1P�s2�*'i~���mӮ��R/�Q,*f-���D���bN�\��}73e�����U򢙉����8�zt�dc��# X��;�a�Qn��2<���і!��]3�nЏ��2��#F�YTf�N��C�(	��-S��j9W�٫>-tPhd9j����)U\�pz�Ћ��obMq=�g�]���[)��}`�+u�u�c����l�4m~��sN=	�8.�_2Y6;���>T y�U�P9��r�\z�����dA��+�å�v
����g�L�����z<Z���B��e��*�:uF�� W')/@���r���*�]��#�Z^��_մUmj lz�9�xt]�d��-Ҳ#�{6��������5&��ٚ��q�����X���m@u3���w��c�%s6��8�p�� $0]5�7�u�pK]�ض$�=z���g�1��� {9	hTʖ�����S��tr�#�25y����#��m˽M��r�6�Yd��	���}�	RU�R�Y({���ۈ�|��z��L��Ҫ�6~^��ڡ�n$�ۭ��Omm�w�Q�,��`��(ᡉ�f�<.Aы 7"���60"���ѕNr'B�~��њ�6i1o�&�O��x(�T�������LH�N�nGf�pfݱ5�I�z���-����M�!<.e�=om��L�$�!dEJ9�V��$c�z�su �'�!��$�B�̡��o��7<s�n���*M�c�&��_��Mc{ؐ��������ڢ�oY_�t�v,l� �p@徏U�n3R
�tR	~R7�}i�\[�W���,����)�B����a#�� Z*����tc�o����E�K�q�
U~4�����u�f�g�˹����*�U��������煦쮗\��B�X��鸤�q;.����PD�{�����ֵ�BJ-,�>��(�A�{��>[�L�L��5�đ�����$Q9P���k���x�
A߾��="ׁ�z��KDՐ�
�a��r������"lA��8�8�G�ܸ�l�p����� V�lj	�(���Q���ȓ�Er* ��r6$�Q���<w��8҄�F[`��d�]P�Bb�����O����PP����}p�4���x�_E`.�a�����<?v'+�@�v��������r�
�;�[XBoP�rհ'}bs����۷-sܐZh���o���!�Z3'��3j�V��^F��B�qW�Q�o3ĦY:��
��^���,iRڙ]EY#��R�u����Jq�7�:��"��Uؠ�F�+mT
|RHt�=��#w��Y��qn7h4v��b8���K<����;#a&�ŦZ�{BJ�-�l� ���#���g�����8$�C��v��6%�\�;��LrDɽC@��C͎�Uo�s5���׍�^��5���N#ч�s�(�k�^+���wi�FmZ-��J5��k�yQ��=�$p5��V����%-K+ϻ�$��Ε����e�c��P����A,�!�:gn�"P���-�Ʀ���TxmLJ���K��0Z�J��}	��V�S���/�����m+��a����dG���)W�C��A��K������[�:��w����,7�^���76���qz����r'�ZJ�U�C8M���i�썚�Rځr�TE\���n2A|�^Zm��a���x]�EC,��S�oM���q�bFע(�da���^;k�iblm�!�{:��OXxdhpǴN �=b®	/
�nrR��ǅ٪N��V<����ƒ.���<j��j��&,(��ڊ��񊪤���4~� )�I۽t�=��&��,v|j�j㉚���8��\d�!�KE�v�	K�EU/P%�V<Z�6��؋o����{w�u��LyKq��� ��@�y�RD���1p߿{�Xm�;	'1V8��֖�8���)pMg���6B��"0GƱ"<;av����vS�����@��Dw5��*,���{V~vq	$�1���v������H�l����r5��^p|أ��<�����.3����*�6,��s���1�9�,���Ч���G�S�Jph<��*��Hl�Dz�y��^�˩�\sǅm���4f6���G���h:qB�﷐�Ѐ��Ķ����8���%�}��6�����I�r��h� ��}L�𣟏��a��Fѽ���M��y�8�RBz.���S�ٗ���|#���b~pe�m�P�B=�P�I7j}�U��JQ��&\`\��W%w�S��c�W��_%�$H�\3zBb���=����q�P����:C4�q��Jr�'����W+��
v[�h�J����
����RV�����u�ދvK=�dl��ݴ׭r�� ��%F<�ǋ=�oh'�p�v���=A\îv*^'!G�@9�zdL���px}N";wx�Z�ps~0�x(8��njt�|"ճ�d�3��^:���[���w�>_��Л�~ٲ�Ie���� Ϊţ����*0#!҂H���W���!L1��`5��t/���q�f5���Y/�|�n��i�*�U=\ȑ>��;��X���΍>��d/��5��q	���}��8e8�B�f^d{�h1i��ѻF�Y�G��c)�/9W��\��EuA-�'Œs��X�B�S���U9��i��[�S����8�K>��^��yy�����.�͙^�����X�6c�Ub�I\�Nv��Nٹ�n����������]a��L$��P5��|���-xG�6I-�-u�YF4�Ss��]m�vVy�Y/�A;��lv�(FT������,J�*<�*��z��6�QS�h�:����t����r'�)�ؓDk�#G�z��9�e���Z�X�]�ƹT;�:v�7�p6�ݡ�ΏA��ٲl��vhO��V���6�d������hd��h��p�0�WdǴ���:�+�&&��Mݔo��9��~V4=�J�M�Y4?b�lu;ђ0QD|h���MF�ԝ�wKjPg�qn��[5;��&�#U����r<F��I2Q8�81p,]o`�ڄ�y9��a���B��ocw
�O>R�����6��v&Ǥ�j+�=S�M�U@
�&]ͻ6�O�,�e(���b���I��f�ߜ���7��2U��98����-�?Ԯ�OZP	b�Ju�Pwe)JM޸�P45|�m݁4 ��k�nnO7)��:�U�3�b�B�` ��.�h��*Eq�Z��<���0�x��1M��Fu�
y���c{�e�@Sz8I7����'��x���Ŋv��������v"l8��Q	�
QvV��c���`l��X0��f�l����I?Z%bk�j�ͥ\!���������A�����á�����.ݍͅ�2��0�t�-���]"�����6�}C�,X�q��^��xҜ����e{w\�W<mn��x�l&��������w�R��h�D���e��G�r�	��"tOvx��=���\p��Qo�ٙ�����@K]��útwM��A�ә48g�8�U�f�8���]۽,�@9���wi%W�\B�{��Q�ᆏ'�g�l�̐x��f�7�}(�%aX�a���]Y�ofZL�A޳���9ԛ)j�>����xD�B������
VgN<�%Y�L`�{]�*HҤ0 ��o�\�&s�n�Λ��\S��	�h&�遤�H�ǈ":�9KM☽|�|�Js{���3�lڌ������{��oq4�/�6��
�]_�Ȩ"�ڃ���z	���{bӑ���kس�����<�����Gtj�nl��VȥB�9M������<��|t
�������C-��t%�I���U���� c�}���8�F���T�oB�#�|��o��N���2�պ��� ⫌�mU�_tG˔&�ա:Y��.�)/�}ޜ����5�}�����F�$���ŘJ�]K�Ձ{�H�}�8��A/�v�ΏD-6�0���2ۆV��O'��=�v��ȅ�KKs��"���;�^3▎!҇q��"ް����ϗ�y���V]����c����Df<d
cdwF2�/5�a{������]���/���f�wpS�v��7Cuc��^�YkXE�ē?*�����`�%5�pk��
��z!fYl�5��X��ɇy��Eg7Bi�6(��5���R#�7���z�@d3T�C����>����b�ⶻ�E�1tj�o�,���o���n):�7�8���ZuݶQ�t	EM�:I><�$���������j�ƥ�~\Z�)x�:�6��0�ƓO�>{Ld�☘�{����Mr�>`0��3� ��}3��؞o��X��6��
�;��4���q6Ao��<���D���jm}���IZ�`@K�$����ϙ�h�6��v��F�1KE��jm��Ү�.)�� �܀ng�غ�6�f*���4n������#�I�C5�PF���0%ʿXxJ�N6�%eg�dI� ������Bl���T�<�ۊ'����=rw{��SBY�{v�͓�C���~�T?i�F?K@j���ч�?\��&{��T~���`��O�����r`p���̴x���]a�!R�;	�]/�*�_��6��� BX�h��%���(;W��MM\ι[�9m{��#�4���P���ј�ѭ���7��K��:�|ŅZ�_n�z ��.'�h�Q\���{`���4�Nu�����#���ۄ��Ʀ�vG���n%��vٝ��lـ�Fz {q��WmK[b�K�>8�BP���� �ډn�@�q�H���Zz J����x;�Y�4�ZoL�(q�-q<��Jr��=(
I[���,�ģ�qݘ�.lj�k;�_c�Gi}��\Hg$�.���~_��&7���sk�N��%{�t'�A�*߸m=^��j7KY���:٬_o��	�'w����ҟ���2z;��X2m���r�8��˳z�͆V��Bz�� �Ʀ�6zm����;�(�<�'+�ካ"�2*zRB��N�����̹8��c��{�2,���lә�(�B� m����Jrd�z�J\�^p�\W��w/Ȏz�F�'������F���T���(w���˩��u�pb�A�F��S���͝9�;7�� |���vK���W�V��S�I��F��;�<��O����C9���B��vA�\o�CrAo�&���w���3$,��5�!�`�*�x����i݃��Q��HN��/$�:��]<%�,5T�؛r��LW����S�U��+q�M��M� �b��q����8����!�ŋ�Mf���E�&H�<��X��q ��F�Q���� G{����o&�!j�n���;�>F�9�u<���X��}������� ���]��Z÷"�6��fl�-�L�d�N�1X�� 9���DJq��/Em��'&b]��1C� 6�u5�T˜a�]�*�Ǟ��I����Vg�";��|�١4�_=T�AwU7Ǎ����~����*��"����٢Yv�/�a�A-��-З�`��2Q����q-�m�cx��a0nG���;���g�
��T�f��|�Y�m{�)�<e[�ǎgÓ�Jh9Z(���f���{�����s��~r'eZ�R����s6�׸�B�n���)}�k����z��s�Dө9�'<��3����X���/�6�������ğp�fNt��(�E��0���}x���sV,z���G9��xz�y ��z��xx>o�r&Gӵ|�Pu�V�N��&�$<���\L(n���#��X��0?Anz<G���緋��Xp�Bz��M�A�����PVC�u�J�F��ƽ���)�L��,ݡ,�}����R�h9A[���K]ߋ�}7`[^�w�-xY��G	̴��Z �3��1��)�����?;��%�͑ɺ([��)���.��1uڹ�eoo�W�P�V&�AG���(��M��/k.$� úA�UU�i�j�r��3	� �3�c��7�v���n?T�a>�7ؽnl���Z=Ђ1U��E�o.�YQUj���&x�N<�l�fZ��]�.���.�q�[}��n#�:���-�P��?Hv���	ou���~R�ຊHP69E��<W��1m0k���&��-[�Ҭ���Bw9������w����6��7-q���f
M�;:A��8-\?
�g#/A�Ё_��10� Vۺ8�����}�$�$�l�y??nU_��579k���al�	RC�ʕm���#����m=AKx^�}�֙�
x���2S2w-��T���ޡ�aP��t�O��AY����U�S��-�V�Iw�q]��O�( =���t�2w��Z���6fd���Ԩ�Ls���*�lѩ����k�_��w�*͖��j�$UTޕ#��u�����Aެž3ʒ�pE@Ǜ��T����޾)Y�"�<�n5��F�2u	��WC��<�r]@�	*�x���-�_&�[~�q��� ���ɪ�o��<�����)_��?�ޣZ�@_~��0�q��`�1��ᑅ"t͠� 9��������X�뵮BҮ�jn>}���޻ʢq�s�N��i������Y�)�0��P8��33ς@�����O����_�aۂ:����|�� q́D�����u�����)	��S1�֜D����{8���\j觬Ʀ W�>�:�Z�_���q̺�C���.ڢeڋ�����M�����or@����U>o �i}�iV�����y���|��-�Y�Pg⋻y���?g3�� {�o�=��G�怇`.>��9�^zd�g�9��cV+� �S���k����;�yG���>\�����g�BxT?�.����s�a��}���{�&j�'��z�|�����n�$]�3B�+WV�Z��E��������X�C�e�y�C_lBY���U^j P�/���,׭ͷ��������J�wh_��ߗg>>]��(p�V��U��k,��eq�# ݫ.�B���k}	�y�g.-|?	v��91��)鰸94x�}f_O@�>���`m�S8��g��W�U=�9 ����~�#܅+((�}�( z	d���3EH_h��T�������/S�_��RqcT{���n����6���"��/h�K�#�=E�-x�EЗ�z���"�q/RĴ%���s�>|[-���S��a�)�YW/��Z�z�����/)�3�~�azi�/Q���{�W���*���SK�������������}Ϛ�A�F�I��^>)��b�/QT��G2�3�(j��0�x�ї�t�h��˳�d��"G�k8 M���.3\/_���/e��M��e�v�ue�K׵%�{��}/���˲��s�柏\��@a/��*��˲4��T�'*�py���GV���@���Z��(.����h��f�q|O�^.���W/P4\myI�<�.�+/s9�gس����>��z�� ?��?1���
`?�ՒT?���8~�w!�}Z��� �Lq���R{����z/�X�%^^ֻ���\���lO/S\-�ZS��^�늶Pt��]�#]my��+H�K�'�p^ֻ�z�?��
��Ji/�]�����])
��z�K�e��5�^���7��w�(>�����C_�� �T���w�e�~�w�(��<���E���D�/P��ap/�]��������݋w���7�b/c �ً���Q���ŀ�G^���A}�b�X}��.�L��&�}���S1V�|=7����������i�P�>$@���?~�M�Qs�+��}�I�6�?�� $��<��n<k>�g*����8T'I-u�B�գ�Δ�-U�&08����Э��I��*h4��ǨY��_t(8�P*��Z�]15�Ym�z����K���ӂ�����x������wį~�z|�J�����2yz}`W�QCV��~�s�/���X��9�{rT����V~�=�͋}\}�����!�����jL+{�?����}��}�g��
���f|�T��:���P��YW�.����yG�KZ}W��]x�a��� �e]���jc���?��7��n��Nz�2ޓ��[�ZG��"� ^A?s�(��=���_��_�o��hu>`�"�-��9�OM�^w�y_jݗ^�N���O�<�5@b�u0�e��d�H����{"��W�}��J�GN v�9����دk�t�3P����q֕�U��uez�ܧM��x�}�a���۩��l���C��縐�O�bi����ꉯbУ���>ף~\W~�2�ֺ�xFW^s��r�/��#�/k�?�f���6�^�gW[}X��[���	��z5��OW[�7k��=?����+�/@]��F_��^���0���~~�2~���5�`}���Sb�[����*�{A�����%���\l0��p:*k���x��|��A_~�ׁV�~�V_������*��W`v>�K2|���[�ֵ�]F��7~mN�:m����6���}��$��o�t�O�V�վm+7�5�%,��خ���?4�/����C�ܰ&�X>o��Ո�M���(�������v�ٍn�1m��^/{�8��4&W����lW::?���\qro���������&#��
1!���(�;�����5?��"����%�n���Pp�#��h�t��3�K���M�O{71���1�@f���#��+Ö��3�SX;�ݘ9��4��s(,�# � !���|����o<�~\p�8���/�m�M�a&��D�я����3�,3�J	�DZ�5k=GI���mn���E�b��1V)1�91�٨S������o	qC8`L���n�M��!�
��19�11��;���O�%`XL��,.�9�̴I�Y��-	�~!�N�}��ǁ���(	�#�R��.Wi���x��P���*�e�?̬BUsX�9��Ǉ��r�u�U*���a�ѽv_�Z��p-�]n{u� �v�Ǩ8w7̇�^7����Ặ��{����8t���x�Zt�ֺ>*~t�İ��-�4l�a
��0�ٞ&|@��06�M)�o����<�f���^�(�F�+�a\�����WG	J&���v�1)N�N��m%`J�b�R��VK����I�8���)�
L��MƠu�Lu�/b"C�/��B��0	��p�"���]�SG���#yw�)_�0�8��$"���y�M��1a~�;�O�Y0�xUoXM���s84�4�7ph���c�b��*m �E��q�h]
�v�2%I����#K$�,v6`�N[�Z�G-֞�2L�@8{���ad��%cu����ꣲo��M�0Eő8�Elm�9�����$-#W�ub�I>O��ax��d"`t�Z�Y�kt�g��Q������lz<�8��;�:��5M��
��l�d��{x�߾����=�?c�d1��~c^�������0��\`Jl�[
��&F�i:{���; y@�e��`-{˥��6j��鱰[���1>S��Z2�2��bEԄH?%8��X����O%0�'e�k0r'N<eA��
��"8Ae���Ab�<�ndwWL�t&�]w�e��4�0@{k��F�la[O �(�كD�s�{�U�x�7K��	g����DwV6�����;�cs|�-�4n��[�.e��`�쪴�p
��!� �U呬+ $�t��X�y�5c[���\B��h	�?&JKaj�2u�z��X�LE��	>���l͵L����^g����`�۶b�����\�P��3�����`J�M��C|l��9x��R;�8"Ï���_�S/խ�;��)�W�(Sk���d�B�s����i��Zӗ���b)c�r�rVaa�dRi\���'���rh�Tw'�w�F��G̠�r���j��?Ĕ�'��"��)��lt��-rcT�I�{���!��3����	g�;g6d:E��l���=�R�y�>��=����HO��)3����ƅ��hqف��8��o�.a�K��unO��6Z��*����N�چx ����_��Aku'm���\�Zj�H�ґJ,g�TZ�n<(=~�7p�[qkLdW�}�I#n��0���&JLoS zp���3y e�QCK��`|����S�?A�-�ktP��e�@�P������vf�`�6�Vb2txK,7>�Wl�i��f�F0�6�Mv�(v`�po@C��wh������R��죌rD��>�!��� ����a�Y�X�'�m�aĲ567��fκo~�q�מ>�2q�G)-԰��%��Q�8e8P���0�M8	�����̛�h< ?��7by��l��gc���F1���Fߪ��:'g�5����
[Q&&��ݓ3��`�Z{�����صvS!s�b�m����� ��]�:���{������XM뜾�w=�v�\h�h�lݹ�P_O��?�S�j�-��jw�
�];=��C�_���jLkٴˁuwXy��I�d��o��q��x���^�kqxf��텱�/w�� �2�I�/�Ǵ�.0�E�]�t�@�:�fk#�lN�i��#�s� �U|�i�[��q����sv��3�;	�����ZCZ"����Z����װAƝI�s#X�<BX��'ϯ�o3u?���ʹ{<p��F!!(b��ņ�P[��kS��Z8�#���~�a������{��8��,����
*^f�hՋee�u���Bc�H�~���T��5Z��	ʘ�����J�^%X5)_����[�[2qGHyB��AG�q#0[[te"�?�vJ�K1����(?�}g&�-w�u8��6]����xBc��J$�ST�e��__�|.�3���ܞj����l��/x훭�8^a���f7h}��k$
P�I�Y1�rģr�f\��u	���K3ޥ��U�\#R�������P(��$�~���27w%� 4c2�`  �N�%<�W/0��d,�C���jG�Og�@������������
0����z��}���؟)<�hǟ(�!�����\��k���A���A�j�/,�D�>?ɘ�?�z:�|}��>_�3���)b��&��T�*�1v�/�h4F����<@��:�����=븬�`xw�S,M������?�X�;���XR����x|ˣ�e�z��Gg�Df�� �=) �'���	�����x����p���Du}���}�G��8����H�߯����m�m��|w/CIV�9��� G�O??Y���ŗ� W�|s��WW���9.?�8.~r!<�S$��_1�����T"��'�9�t�V^l���Ivm��c��p��ʨ��+{c$��,6_i��1 /��N`��3��y	������}Q'���G��X5j��~�O����]��I��C�Q�
V�
����O@�?�|$�Q�ӰKV�W>~%	=�>b�/q��D�}_T~��[Z����%�x����~л@u��2�f�W��3f�ʹz��c�90�1&��5&�X����iqҺ�j�pFm�˚�˘��ff3k�?�2Z���at�A&>c�!&~���L@�[1�[���+OB�8�e ��k[��rPX�ZΏ�(a� �$���6��3a���3��Ζl3I�b��1g��5�9�"2J�����ΙT��!�4���r9�3`1�l70}�M���0f�3w��2�������̒�֤�������Ef���}f��df���eI,�	
c��� 
b�+iBl�V��&sZv 1p]����ւD��z�mE�:����K�)��_�tĞ[ǚ=�>[Ē>�A�+)�N$�N��
�LBVT�wOf�����^��"���	�J,^�=�nYZ�q�q̠�S6sB��Y~�E�����1��g��T5綪;�����ZNM�E��L��;;�j/\	�Lw�Za�0�7x;��n�J6�,�C��}Fw`�
��krx�լ�󲧕�|�5FC�e�-HW3����0����>Mhʟ3C�0���2N���3��o��YT�C�y�h��s��&��,�fAЬ �A z㏂�����ף����l˭�Ŏ����XN��Ja���׬��C/Ls;������vA*/̝����%w'�V:{��cvh>-��x��ʏ��{Ň��Ѳ�ZĪ��7}~v�mH���$/(��.�^�ɫL�S�hl)�O(p���=�C�v?H+2c	0&�FC~eF�w�Ñ�!n�&�^"�,���Q^N�T�qFnڴf��|����Hu~��f7[y�f�ò�4e����2'*���[G6��P��zPZ���}�Lmipz��V9&�*KU�cS�n���SU7�C�?�q\�spQ���Uo�E�UE��u>�;j�9�v
�`��vnօs����-�k�k3��nRz����3�{��b.�z<����x�Q���yps9����,�j������-6�.;h;kB�Ѽ������yW���3�k���7����� ���UBx��=Η#��!D_N�~�+a�>��y|�Z��n��+9R����F	��E�ݱ7��$��bJ��Ki:
�Hn��F��̼2��r�'ܖ���t�$p�e$���V�`�J���ʍ����?{&�ݺ`C���p����}�D�
 ���D�B�d/9�ΫC�8Pa;z��^]:a�RB�:x�XE��Mu/\���j&\K�٩�M���7�OLF�U�M��\<Y�n� y�n`��J�9�{�{��6����Y�c�}s��p��C��<|��ڧ�D8����/��W��ק����%����CT���?������$I*��1��H$��D���f	�Cv@�k`>r���|(w���l�ʒ�훓Qצ�;�4iL?tN��b��{�ԭ�~h<:i��,^�z�I�"�K���2�#+3�<h4DH!z��T��17N���b�{�Gy��q�.��r�-oEˋ�Ip�1�#����ȉ��:&�[�=�ݥQ�4!�˵N'��;w�D*;.�������F�L�<c6�<`�lW�\+�Y�p��s���0�ȁ���̽T�b��_v��d�oVɻB#Tk�OR���I�w�����N����-�(O����So7i�c��~�n쫪����`��WdFWQ�]m:�#~T��<�ը��\k��IU�9�a����E=>���i�.�.�T؀�9��h�&Cv��Fa�^w~;�er5�N��a]�4�5�ww�]��Uܵ�]�^���ʻ�y�v}޻^�h}T��!�����ٟ�^̆$�r�K���U����{�f�$$��iD
�秛.�N�n���v#RJ���n�tIb�{�l�$MܷG&��a����7��������=DYX�����=D���;���~Q����܍Ԁ�d���/�Qcy�f�#S�6�y�X�Q���tLz�B��>F[�����6\}DObx�'�l9QI� �{��M�O"��#>�/i;RJl3��ј�拡��x/����Ym_�3��o�'.�v+��o/� ���۱��;I*�(�HL�m4h����7��:���N����Z��a�<�t��;�l�݆�`W��6�8l��=S�v�΅����v\��y��%q�H����)[Q3u��|���t��?�L�{g�a}��Xb6Ƅ�p�Y��Yg��)�z�g<�S�=�ZV��Ga<3?�:��*5BT?Sμ�`�P����0El�����ݫ�t�|�h�i���=*^�5���ы�3e��W��'0��_�Zٚ3X6͉�f�L-���L	e����@,.[�Z�k��g͒�D����ۧQ�.>��@�ݏW�<4�b�H��d�jZ��!3vb��<�m��^��:>&sy4�dOÈ=R���ES���m��1.�B��`F�+1oOd�Jʩ�C�_*bo\:�!+�S17�;)���y���uq;�!����x���$����:Y����*4��K6�˔�=_�����?��b�{���e  ���՛��P�ntA!$
P���l	�������j�"yZR��Y��3�զ��o�	C����&	��N��A�/��DF2��Ac4����iQ>��F��a|�[ި�0��m�Iϼ9)��������~yl���ӌ��b��a6�L*��c��tuƳ��o�+׋�� �� ��Y7�aD@e�:v�*XvypS��,�Mf��Κ���x�|��tɃ�ܾ3���}V�)����֪�9��9h�
v�p�p�b�a� �=6MI)fZU-�Vb�	�8�t��j�&��'@��i����I�LI�ժ|ك�ҡJ��� �������ig�����ܞ���9z7ч={��E�bT�wT�$�	��������
q�S�4��b��v�ԛ!}޾A%��n��F�8O��ls�!G�Kʧj���u��*��(|�v�t�,�y�57��D% yВ`>V\o�K;[e�3�+)�O�z�Н�v>_��c�Q����6]�~rWI�B�2�w�r�����zAW\/�.7���5�ݘ��vG�{��^>�f!��4�dKf��Bq? 9�s���p_Lƌ��T_�H����)uTJ��bZ?/����,�ѲFQ�j�=�v0��1�ǟ��D����F>�Ŏ|q6����u�8� A���}x
�"���k�gq�����~F_H�hf��.q�޻� �n�h�l��U2�Ƥw����*q��쭒�<s����I��p&v����N�Cl���N��+%|�a��e��Yr��X��Fͅ��dםS]�y��l;
��'�N-�EK�y�D�p톼�
�ѭ�F�U��0͌��2)� ���k�:�`��C)�ȹ�Łq� ��[�^3wϩ�ր?}���t �� ��~�F�8�GKL�?n�l#�d0�'y�)?]d)�����*������BO6*���Zb�a�������j,��}�nF0�w���j�I��U�;�Ԇ`�rQ��$��`�J�0x���ba�@j�¸�I�#�9h��w���F�P�2 @c.W�n��@C��L�\+\ �6��᰿BP_^�&����v�����}@����jY�ܐ;rj��n#�T4�wV�j�QA�ܣB�����a�.J�W1,8i��T@W��Pw��I�:=%4�H:|Bk�����Ep�����4lq��.�%#���5 �T�½kw��<w��D&ln�^"L;W���HŜN[���gJ�n)��p�`��x`� ���U+�2@Z�ɥ 	v�S���  "Z8�+\91��hSr%��}=j]�v��/`��St��z{f$�9O���f�xu-�DM@6�52�c|
`�"�.L���HL�q.�>֘�d�`��	�=���5~�1n�:��LG��()`�e��L��))S��K�������Hk<s���̌�N�_2�����1Q =��&�4��d{�	K�>�Q4�Cj{����ْ����M/UXH��X�z �\A�&�\��YG�Pi�Rq�PU��+W�KS��Ή;ҹ.;����1ukf��������R���{���S��p�l-�S��͒�z{��k=��]b����zW�!X���{O,� ��5���GY�M?P�Q��}J�F�ݘc�v:�z]���z�K�,�<F!�h�<�W~�] �4�R���@����v�L�+qCk-y$��� 7J�r�N����U���v�5y;����țT��V��z|74mu��=��b��T��1������mƘ���޾�k����8��12�Q䠅?�Ӂ�Q��$&G��2����K�Ɲ�w��(�0��f}�e1�C-���g^=��5��{��5McZ�[ֈ2�F���������� �=Yr�d�L��4We;���0��z�53+���rj֘D�9l��d�t;X��$Kk��gVj�\v\�l8q�1Ӄ�MA-4����'�����|!�����؉�#p���u��ǭ��G�>�+��y3Ku1��&�S���V�(g����� �U��Y8V��C�̧T��1�.`�.7wm��W�]䶵��e	��@2�zޝ�L� ��kd
՗m������� Zڱ���;ێY��jغ"��="qI��jE]�ET�X���Ǐ\u~�F��Wf���Y,�Ă@���'��?�m_��}��-D�Ll�����yL��ə	�-A^�9��zV��@�v��^�"��ŕ�Jm�7j�?�]ҿ}ӘװT����~�o��:^�cG;]�a�H7���C{��} �����~r��X���\��a<K��Ҧ�r��E�z#ɘ\��#rA7��J���.I�5Y�t�M:�ýVm��1������Ob���F�X�Z��#S�s���{�l�)cj,�	Ū@׽F��l7�"�zk)�������L����虍"�PjX�9?�<>�j�f��,�ɗ5�/z�hUG�8����\��w�(0��f �(fp� ��� (��7�\Ԅ�s{P��s']���O�x���#$m:Ey�J���ɑ5&�Y,�G�9k�48pͬ�
����Uj':���FN��2�
9�d/U�>c�~��}ɉ���R;i�ػ<�z�ץh�#n�]3�ޔ�o��ԍE$���J 5��w{�� �Z�[r2��(q����_Հ]m6�����T��(P �j�I��Q��Pd����H��+B�b	z>�\�WM��~:��P��Z�*���C��g��[��n�Z���w:V[�ߩ�I���8�^'����a]�Ixu�+.J�m�4R�#�"�q�t&ae�ę���pepGL\Z����!vkoӇ��،� d����e��.N�bLY�'���hm�l�������y���r*���CG^Xc���E��������l���>+6c�ᙷo"	#���\r}l\ܶ��Yi��几���i��z���>�}q��S7�c��퇖N����]������$E<�o�7cⱸ��pN{咤��'����&��O�?��~>�6�LRކ����n?�aø���vI�>��"���N|h��>������������KAĿ������w��|���Nwں�|��NS�/��x�����a8ǹN�l���7�0i�/Z|��}��/�����{~���c�V���_����sd��=��Ȋ���qz�����g����0u�]^`(��z�Ӆ1 ��9}�����}��Ԝ/`�f'����݂��$�Kq��������/k������Wl�IT^����N�I�
Q��
�+���;G߱��<��i�K_�����a��o8��& �^����cx����"n��l߶�<��3���2�q����%n�6\��P���p��1�Co��_��e��/g�/�a*��/�8�!�_䴾�c�����q[�=h����O�Z���izY�D�-���_��O�2>p�ay���� ���}6A�g{6��gp��B��&	�\�'颿���o���~�K|�~qnѿ�m�_�M��:���̅�2ן���\���wL�C�ye�:{�Eݎ���&�A$@q��Q(���4���� ��m��]xǰw(�^�?��?�dB����4��g��Od�W6������Hb��8���'���`pA�(F#�YMi�,���s_\���٭�_��f�������Wc&Z�]�����ƽ�b��z�$!��������/��p� ���!��~�-���3���B�m���:�7��e�E�~�z0�z�*�mY�K:|{�g �"��� �0m�r��/`z`�����[:�]������Um�mjs;�}��p#'��!�&��7_���|՛��ބ�ŉ��3��#��!��"8�s��W���dy��_;�[��Ηj���"Q.���υ�������v�����7O.e���7>~ܥi��>N<������c��7>*ܷq��~�$vm��͋�-D�%�~�|0�tη#���H����gs����?�5�R4ᘾ0g����y\�q���ǰ������I�c�^�; ��Ω��.��/�+i�:vI���8�]����g��H/�7g�(1�3�te��p��N��x��7?�&����҃x���b��������l�<ۻ��W��;�6��<���.�t�oq��6�#Y��[Mܯa��e<	��� ȿU�������A�w���	ëHa(8�~o+�w���vX���e;ˋ Vx�k������7x�k/^��O��;"OU�/O{oؑ�\��e���?����@~M�K���|���P|c�?�q� q����)��P�k��}o�ݹK_���O���[�㷅%����ט¿�����_��@���-0���_�j}����� Suȵ��f *�ow��g��(�����#_��/���J�Z�U���ь��>�-AVA��(���q��V������蟷D>�$��Z���:�7I���	������e������ �aQ��|�7+�����8�_ϙ�[x��W>���_��;�Vy�V����Q����P����V0~�gC8D�(�c&Y�B=�?Qq߹9_=bz��恒ގ�/������v��	�@�Ίk~y������_�]�a�7@��Y�QzuR!`�i|p[� ^/���"�Չ�=S3��3���o�[?�� �7K��hZ����Y|�u����u}z���tn�/o={����"9����n�ѻ����>{���}�����ҟ�2G�P��+({e2P���@�1���p�U�_�O&��K�)⽀�a����?�Y`{�?L����*&��$�M����{"�@�k,���i�5��x�E����7�"��X�"�H�� �|���3
��L��L'��~�L'�"��L'Ga��`��)!H�5��5��_\#���/�m|z��iN�_2	��L&��Ռ��`�I$
v�X�����JE��Z����T<g��#�.��^S�����s��^�݅�ݍ��/�3����ïm�;��j*�oo�K<�qU�O������b�R���;�x�P��3̆�q���:���˞�g]��"��_�?����O�5����Lb��?�@��}���N����E���|��֓����i�_/����??��}k��>�~�~"�/i���o5�������^��z�[����/��~�7�t�_��[r��&�����x����k��g*��Q��"x��O=����_�~��o5��*����"~?��56�ܒ�_���P�߁�P�9C��^��(��P.���EC���W��=���_�����qp�������Ғ�o�n?��W>��|�R���X�'���Mi֍�_�T�^�y��׹�~�n/->_�+�������/�~�/������i��������k��o�e�;~�d��?8�ï��?S(���w��~����}���Tȕ��Қ��y��Mk����G�P���|�N埰����W����7�ǒ�O�͠�;
y/�Ț�B�C1��_�������m��<cڼY/�������o��ۓ~����l['U�
��f���k�~B_�^��_��M���4L��ũ��#�?�>�]��u��?,3.��ցC鑭O��2��Z�#|h����A"�u�� �|�]�GM�|l�X�[�f�tu�ZL~�	>s?4�p[+��:+���c��h���z�uϳ5p��:���C�����_�U��u�����H��Tޟ-���y���rF,���?4�����gk�Q���P����OݽG���x���=�6�8.>�9�6���E�e�Pzߧ������Y?r�d�?��Z�ڏ�e�γ��
�����o��F�>�nİ�z�0l�HX��
M��	#�%�90.��L\Ĝ�>��I����y܈���)u(��:^����MO��ͣ�$q�d����z��G�/���Z`B��汔��z8Y�ۼ�.�q"��R����󙩿��?����d|=3,��q��wa4�����+y_��<�}���x-��Z6�Tٌ��xfFoW��WU�@^�f�V�x���Z5�o�׎z��?�1�����8�?0:���y���&��l�?ئ��Þ�q�irN������������%�g�9�*�r���?�v��.|���rN�����������s��n[��1��8�5˿zUK�uk�W��-�x������tߺ7K8���;����{��a��p��i����m֖8΀|��쵸�_�o�� o�d�=��R�^y�S�m�q�[���}{�j�u����֙�����ۿ�F�5a^}�?����/����U�yE)�a^Q�+J�WF)�6JA�w�>|,��3�����k��Z��*���j��S��5���)����3���@,����u��¯�ؿ����w�B�*�jP_K���W��{�:���&�̿��D��
�<�o!�����C�����0��!�����&���N^라�;��7�Fp�I���;�����!��_7�~�{�Y�����W�z����F�!$�+��a�0~�"W���X�uP~�B�w$��X��P���P>�3I�#P�B�s�+?�~uQ>������35F�G����k����UR���O>���>�k���(ؿt������?~���~Q�	��u�^*�Tx-��g+��끏��݃�
��V�prpm^�][��D��Q#~���>7�;߭%>WMhC�S_��p�B�!Bf�`0���nn-{�G�"���F�G�� Q.�������ǫ��v��-��]��NM�_��jN��V& }�@��OTp�C������9��b����50$����3��akF�>v7���l1�Ŗ�$0{���b"��>���qi�n-� E�:0�c}h�m��g݃ |���&"6�x�_N��k/|� �Q3��ϗ��BoZ��A,Hg�Iar���6x-���S��D�繙��^��z��ZHᵐ�k!��B
�^Ha��@e�U�ߡ��g�}��(���7`x�[�����
I�,�O^y3���_y�7��e,�������8-.� ~)Q��齁��=��s�?���`�Zxt�%I���1l_��oE����-1}��p����7οUC_����%�;����@8ԇ:���I~���^����JS}�X�^Dnc��/�1a80����,0qQ�ٽ�BD>��V���.����Q����~P�Cթ�f_������5����������`/�ةm��g�ך���S�C �����-3��U^��+���%~Ve����K�篦��.��^��5��֭��}�VbQ��Ǔ�c�Հ�����I6��^� 